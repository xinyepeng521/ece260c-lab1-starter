module asqrt_top (clk,
    ready,
    reset,
    valid,
    queries,
    results);
 input clk;
 input ready;
 input reset;
 output valid;
 input [127:0] queries;
 output [127:0] results;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire net24;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire net23;
 wire net22;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire net21;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire net20;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire net14;
 wire _0151_;
 wire net13;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire net12;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire net11;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire net10;
 wire _0169_;
 wire _0170_;
 wire net9;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire _0183_;
 wire _0184_;
 wire net4;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire net3;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire net2;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire net63;
 wire _0204_;
 wire net266;
 wire net243;
 wire _0207_;
 wire _0208_;
 wire net62;
 wire net55;
 wire net53;
 wire net242;
 wire _0213_;
 wire _0214_;
 wire net275;
 wire net59;
 wire _0217_;
 wire _0218_;
 wire net274;
 wire net273;
 wire _0221_;
 wire _0222_;
 wire net260;
 wire net58;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire net268;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire net276;
 wire net261;
 wire net272;
 wire net267;
 wire _0236_;
 wire _0237_;
 wire net269;
 wire _0239_;
 wire net265;
 wire _0241_;
 wire net264;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire net262;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire net259;
 wire net258;
 wire _0301_;
 wire net257;
 wire net256;
 wire _0304_;
 wire net255;
 wire net57;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire net254;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire net253;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire net263;
 wire _0381_;
 wire _0382_;
 wire net252;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire net251;
 wire net250;
 wire _0389_;
 wire net249;
 wire net248;
 wire _0392_;
 wire net247;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire net246;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0465_;
 wire _0466_;
 wire _0468_;
 wire _0469_;
 wire _0472_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire net34;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire net33;
 wire _0568_;
 wire _0569_;
 wire net32;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire net31;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire net30;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire clknet_0_clk;
 wire net1;
 wire \genblk1[0].pipe.counter[0] ;
 wire \genblk1[0].pipe.counter[1] ;
 wire \genblk1[0].pipe.counter[2] ;
 wire \genblk1[0].pipe.counter[3] ;
 wire \genblk1[0].pipe.counter[4] ;
 wire \genblk1[0].pipe.eps[0][24] ;
 wire \genblk1[0].pipe.eps[0][25] ;
 wire \genblk1[0].pipe.eps[0][26] ;
 wire \genblk1[0].pipe.eps[0][27] ;
 wire \genblk1[0].pipe.eps[0][28] ;
 wire \genblk1[0].pipe.eps[0][29] ;
 wire \genblk1[0].pipe.eps[0][30] ;
 wire \genblk1[0].pipe.eps[0][31] ;
 wire \genblk1[0].pipe.state[0] ;
 wire \genblk1[0].pipe.state[1] ;
 wire \genblk1[0].pipe.valid ;
 wire \genblk1[1].pipe.counter[0] ;
 wire \genblk1[1].pipe.counter[1] ;
 wire \genblk1[1].pipe.counter[2] ;
 wire \genblk1[1].pipe.counter[3] ;
 wire \genblk1[1].pipe.counter[4] ;
 wire \genblk1[1].pipe.eps[0][24] ;
 wire \genblk1[1].pipe.eps[0][25] ;
 wire \genblk1[1].pipe.eps[0][26] ;
 wire \genblk1[1].pipe.eps[0][27] ;
 wire \genblk1[1].pipe.eps[0][28] ;
 wire \genblk1[1].pipe.eps[0][29] ;
 wire \genblk1[1].pipe.eps[0][30] ;
 wire \genblk1[1].pipe.eps[0][31] ;
 wire \genblk1[1].pipe.state[0] ;
 wire \genblk1[1].pipe.state[1] ;
 wire \genblk1[1].pipe.valid ;
 wire \genblk1[2].pipe.counter[0] ;
 wire \genblk1[2].pipe.counter[1] ;
 wire \genblk1[2].pipe.counter[2] ;
 wire \genblk1[2].pipe.counter[3] ;
 wire \genblk1[2].pipe.counter[4] ;
 wire \genblk1[2].pipe.eps[0][24] ;
 wire \genblk1[2].pipe.eps[0][25] ;
 wire \genblk1[2].pipe.eps[0][26] ;
 wire \genblk1[2].pipe.eps[0][27] ;
 wire \genblk1[2].pipe.eps[0][28] ;
 wire \genblk1[2].pipe.eps[0][29] ;
 wire \genblk1[2].pipe.eps[0][30] ;
 wire \genblk1[2].pipe.eps[0][31] ;
 wire \genblk1[2].pipe.state[0] ;
 wire \genblk1[2].pipe.state[1] ;
 wire \genblk1[2].pipe.valid ;
 wire \genblk1[3].pipe.counter[0] ;
 wire \genblk1[3].pipe.counter[1] ;
 wire \genblk1[3].pipe.counter[2] ;
 wire \genblk1[3].pipe.counter[3] ;
 wire \genblk1[3].pipe.counter[4] ;
 wire \genblk1[3].pipe.eps[0][24] ;
 wire \genblk1[3].pipe.eps[0][25] ;
 wire \genblk1[3].pipe.eps[0][26] ;
 wire \genblk1[3].pipe.eps[0][27] ;
 wire \genblk1[3].pipe.eps[0][28] ;
 wire \genblk1[3].pipe.eps[0][29] ;
 wire \genblk1[3].pipe.eps[0][30] ;
 wire \genblk1[3].pipe.eps[0][31] ;
 wire \genblk1[3].pipe.state[0] ;
 wire \genblk1[3].pipe.state[1] ;
 wire \genblk1[3].pipe.valid ;
 wire net164;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net54;
 wire net60;
 wire net241;
 wire net56;
 wire net52;
 wire net61;
 wire net64;
 wire net244;
 wire net245;
 wire net270;
 wire net271;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net277;
 wire net278;
 wire net279;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_tielo _1226__12 (.L_LO(net63));
 sg13g2_inv_2 _0648_ (.Y(_0204_),
    .A(net276));
 sg13g2_buf_4 place266 (.X(net266),
    .A(\genblk1[0].pipe.eps[0][29] ));
 sg13g2_buf_4 place243 (.X(net243),
    .A(_0574_));
 sg13g2_a21o_1 _0651_ (.A2(_0204_),
    .A1(\genblk1[3].pipe.state[0] ),
    .B1(net270),
    .X(_0006_));
 sg13g2_a21o_1 _0652_ (.A2(\genblk1[0].pipe.state[0] ),
    .A1(_0204_),
    .B1(net270),
    .X(_0000_));
 sg13g2_inv_1 _0653_ (.Y(_0207_),
    .A(\genblk1[2].pipe.state[1] ));
 sg13g2_nand2_2 _0654_ (.Y(_0208_),
    .A(net276),
    .B(\genblk1[2].pipe.state[0] ));
 sg13g2_tielo _1225__11 (.L_LO(net62));
 sg13g2_tielo _1218__4 (.L_LO(net55));
 sg13g2_tielo _1216__2 (.L_LO(net53));
 sg13g2_buf_4 place242 (.X(net242),
    .A(_0128_));
 sg13g2_a21oi_1 _0659_ (.A1(_0207_),
    .A2(_0208_),
    .Y(_0005_),
    .B1(net273));
 sg13g2_inv_1 _0660_ (.Y(_0213_),
    .A(\genblk1[0].pipe.state[1] ));
 sg13g2_nand2_2 _0661_ (.Y(_0214_),
    .A(net33),
    .B(\genblk1[0].pipe.state[0] ));
 sg13g2_buf_4 place275 (.X(net275),
    .A(net270));
 sg13g2_tielo _1222__8 (.L_LO(net59));
 sg13g2_a21oi_1 _0664_ (.A1(_0213_),
    .A2(_0214_),
    .Y(_0001_),
    .B1(net34));
 sg13g2_a21o_1 _0665_ (.A2(\genblk1[2].pipe.state[0] ),
    .A1(_0204_),
    .B1(net273),
    .X(_0004_));
 sg13g2_inv_1 _0666_ (.Y(_0217_),
    .A(\genblk1[1].pipe.state[1] ));
 sg13g2_nand2_2 _0667_ (.Y(_0218_),
    .A(net276),
    .B(\genblk1[1].pipe.state[0] ));
 sg13g2_buf_4 place274 (.X(net274),
    .A(net273));
 sg13g2_buf_4 place273 (.X(net273),
    .A(net270));
 sg13g2_a21oi_1 _0670_ (.A1(_0217_),
    .A2(_0218_),
    .Y(_0003_),
    .B1(net275));
 sg13g2_inv_1 _0671_ (.Y(_0221_),
    .A(\genblk1[3].pipe.state[1] ));
 sg13g2_nand2_2 _0672_ (.Y(_0222_),
    .A(\genblk1[3].pipe.state[0] ),
    .B(net276));
 sg13g2_buf_4 place260 (.X(net260),
    .A(\genblk1[1].pipe.eps[0][30] ));
 sg13g2_tielo _1221__7 (.L_LO(net58));
 sg13g2_a21oi_1 _0675_ (.A1(_0221_),
    .A2(_0222_),
    .Y(_0007_),
    .B1(net271));
 sg13g2_a21o_1 _0676_ (.A2(\genblk1[1].pipe.state[0] ),
    .A1(_0204_),
    .B1(net273),
    .X(_0002_));
 sg13g2_nor3_1 _0677_ (.A(\genblk1[0].pipe.counter[1] ),
    .B(\genblk1[0].pipe.counter[0] ),
    .C(_0017_),
    .Y(_0225_));
 sg13g2_nor2b_2 _0678_ (.A(\genblk1[0].pipe.counter[2] ),
    .B_N(_0225_),
    .Y(_0226_));
 sg13g2_and2_1 _0679_ (.A(net33),
    .B(\genblk1[0].pipe.state[0] ),
    .X(_0227_));
 sg13g2_buf_4 place268 (.X(net268),
    .A(net34));
 sg13g2_nor2_2 _0681_ (.A(net34),
    .B(_0227_),
    .Y(_0229_));
 sg13g2_nor2_2 _0682_ (.A(\genblk1[0].pipe.counter[3] ),
    .B(\genblk1[0].pipe.counter[4] ),
    .Y(_0230_));
 sg13g2_nand3_1 _0683_ (.B(_0229_),
    .C(_0230_),
    .A(_0226_),
    .Y(_0231_));
 sg13g2_buf_4 place276 (.X(net276),
    .A(net33));
 sg13g2_buf_4 place261 (.X(net261),
    .A(net260));
 sg13g2_buf_4 place272 (.X(net272),
    .A(net271));
 sg13g2_buf_2 place267 (.A(\genblk1[0].pipe.eps[0][28] ),
    .X(net267));
 sg13g2_nor2_1 _0688_ (.A(net267),
    .B(net266),
    .Y(_0236_));
 sg13g2_o21ai_1 _0689_ (.B1(_0236_),
    .Y(_0237_),
    .A1(\genblk1[0].pipe.eps[0][31] ),
    .A2(_0011_));
 sg13g2_buf_4 place269 (.X(net269),
    .A(net34));
 sg13g2_mux2_1 _0691_ (.A0(_0237_),
    .A1(\genblk1[0].pipe.eps[0][31] ),
    .S(net265),
    .X(_0239_));
 sg13g2_buf_4 place265 (.X(net265),
    .A(\genblk1[0].pipe.eps[0][30] ));
 sg13g2_nor3_2 _0693_ (.A(\genblk1[0].pipe.eps[0][25] ),
    .B(\genblk1[0].pipe.eps[0][24] ),
    .C(\genblk1[0].pipe.eps[0][26] ),
    .Y(_0241_));
 sg13g2_buf_4 place264 (.X(net264),
    .A(net263));
 sg13g2_o21ai_1 _0695_ (.B1(\genblk1[0].pipe.eps[0][27] ),
    .Y(_0243_),
    .A1(_0239_),
    .A2(_0241_));
 sg13g2_o21ai_1 _0696_ (.B1(_0008_),
    .Y(_0244_),
    .A1(_0239_),
    .A2(_0241_));
 sg13g2_inv_1 _0697_ (.Y(_0245_),
    .A(_0013_));
 sg13g2_mux2_1 _0698_ (.A0(\genblk1[0].pipe.eps[0][28] ),
    .A1(\genblk1[0].pipe.eps[0][31] ),
    .S(net265),
    .X(_0246_));
 sg13g2_inv_1 _0699_ (.Y(_0247_),
    .A(net266));
 sg13g2_o21ai_1 _0700_ (.B1(_0247_),
    .Y(_0248_),
    .A1(_0245_),
    .A2(_0246_));
 sg13g2_or4_1 _0701_ (.A(\genblk1[0].pipe.eps[0][26] ),
    .B(\genblk1[0].pipe.eps[0][27] ),
    .C(\genblk1[0].pipe.eps[0][28] ),
    .D(\genblk1[0].pipe.eps[0][30] ),
    .X(_0249_));
 sg13g2_nor2_1 _0702_ (.A(net266),
    .B(_0011_),
    .Y(_0250_));
 sg13g2_a21oi_1 _0703_ (.A1(net265),
    .A2(_0013_),
    .Y(_0251_),
    .B1(\genblk1[0].pipe.eps[0][31] ));
 sg13g2_o21ai_1 _0704_ (.B1(_0251_),
    .Y(_0252_),
    .A1(_0249_),
    .A2(_0250_));
 sg13g2_inv_2 _0705_ (.Y(_0253_),
    .A(\genblk1[0].pipe.eps[0][31] ));
 sg13g2_a21oi_1 _0706_ (.A1(_0253_),
    .A2(net265),
    .Y(_0254_),
    .B1(net266));
 sg13g2_nor2_2 _0707_ (.A(\genblk1[0].pipe.eps[0][31] ),
    .B(\genblk1[0].pipe.eps[0][30] ),
    .Y(_0255_));
 sg13g2_nor4_1 _0708_ (.A(\genblk1[0].pipe.eps[0][26] ),
    .B(\genblk1[0].pipe.eps[0][27] ),
    .C(\genblk1[0].pipe.eps[0][28] ),
    .D(_0255_),
    .Y(_0256_));
 sg13g2_a221oi_1 _0709_ (.B2(net267),
    .C1(_0256_),
    .B1(_0254_),
    .A1(_0248_),
    .Y(_0257_),
    .A2(_0252_));
 sg13g2_buf_4 place262 (.X(net262),
    .A(\genblk1[1].pipe.eps[0][29] ));
 sg13g2_inv_1 _0711_ (.Y(_0259_),
    .A(_0011_));
 sg13g2_o21ai_1 _0712_ (.B1(net265),
    .Y(_0260_),
    .A1(net267),
    .A2(net266));
 sg13g2_or3_1 _0713_ (.A(net267),
    .B(net266),
    .C(net265),
    .X(_0261_));
 sg13g2_a21oi_1 _0714_ (.A1(_0260_),
    .A2(_0261_),
    .Y(_0262_),
    .B1(_0253_));
 sg13g2_a21o_1 _0715_ (.A2(_0255_),
    .A1(_0259_),
    .B1(_0262_),
    .X(_0263_));
 sg13g2_nor2_1 _0716_ (.A(_0257_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_mux2_1 _0717_ (.A0(_0243_),
    .A1(_0244_),
    .S(_0264_),
    .X(_0265_));
 sg13g2_nor2b_2 _0718_ (.A(\genblk1[0].pipe.eps[0][27] ),
    .B_N(\genblk1[0].pipe.eps[0][26] ),
    .Y(_0266_));
 sg13g2_or2_1 _0719_ (.X(_0267_),
    .B(_0263_),
    .A(_0257_));
 sg13g2_a22oi_1 _0720_ (.Y(_0268_),
    .B1(_0266_),
    .B2(_0267_),
    .A2(_0241_),
    .A1(_0239_));
 sg13g2_nor2_1 _0721_ (.A(\genblk1[0].pipe.eps[0][26] ),
    .B(\genblk1[0].pipe.eps[0][27] ),
    .Y(_0269_));
 sg13g2_o21ai_1 _0722_ (.B1(_0269_),
    .Y(_0270_),
    .A1(_0257_),
    .A2(_0263_));
 sg13g2_or2_1 _0723_ (.X(_0271_),
    .B(net265),
    .A(\genblk1[0].pipe.eps[0][31] ));
 sg13g2_a21oi_1 _0724_ (.A1(_0236_),
    .A2(_0270_),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_a21o_1 _0725_ (.A2(_0268_),
    .A1(_0265_),
    .B1(_0272_),
    .X(_0273_));
 sg13g2_a21oi_1 _0726_ (.A1(_0265_),
    .A2(_0268_),
    .Y(_0274_),
    .B1(_0259_));
 sg13g2_inv_1 _0727_ (.Y(_0275_),
    .A(_0239_));
 sg13g2_o21ai_1 _0728_ (.B1(_0270_),
    .Y(_0276_),
    .A1(_0267_),
    .A2(_0275_));
 sg13g2_xnor2_1 _0729_ (.Y(_0277_),
    .A(\genblk1[0].pipe.eps[0][28] ),
    .B(_0276_));
 sg13g2_o21ai_1 _0730_ (.B1(_0277_),
    .Y(_0278_),
    .A1(_0271_),
    .A2(_0274_));
 sg13g2_xnor2_1 _0731_ (.Y(_0279_),
    .A(net267),
    .B(net266));
 sg13g2_nand2_1 _0732_ (.Y(_0280_),
    .A(_0239_),
    .B(_0279_));
 sg13g2_o21ai_1 _0733_ (.B1(_0280_),
    .Y(_0281_),
    .A1(_0013_),
    .A2(_0239_));
 sg13g2_inv_1 _0734_ (.Y(_0282_),
    .A(_0008_));
 sg13g2_nor3_1 _0735_ (.A(\genblk1[0].pipe.eps[0][30] ),
    .B(_0282_),
    .C(_0266_),
    .Y(_0283_));
 sg13g2_o21ai_1 _0736_ (.B1(_0253_),
    .Y(_0284_),
    .A1(\genblk1[0].pipe.eps[0][28] ),
    .A2(_0283_));
 sg13g2_nor2_1 _0737_ (.A(\genblk1[0].pipe.eps[0][28] ),
    .B(_0255_),
    .Y(_0285_));
 sg13g2_o21ai_1 _0738_ (.B1(_0285_),
    .Y(_0286_),
    .A1(_0282_),
    .A2(_0266_));
 sg13g2_nand2_2 _0739_ (.Y(_0287_),
    .A(_0284_),
    .B(_0286_));
 sg13g2_nor4_1 _0740_ (.A(net267),
    .B(net266),
    .C(net265),
    .D(_0011_),
    .Y(_0288_));
 sg13g2_or2_1 _0741_ (.X(_0289_),
    .B(_0288_),
    .A(_0262_));
 sg13g2_xor2_1 _0742_ (.B(_0289_),
    .A(_0257_),
    .X(_0290_));
 sg13g2_nand2_1 _0743_ (.Y(_0291_),
    .A(_0287_),
    .B(_0290_));
 sg13g2_nor3_1 _0744_ (.A(_0271_),
    .B(_0287_),
    .C(_0289_),
    .Y(_0292_));
 sg13g2_a21oi_1 _0745_ (.A1(_0287_),
    .A2(_0289_),
    .Y(_0293_),
    .B1(_0257_));
 sg13g2_nor3_1 _0746_ (.A(_0281_),
    .B(_0292_),
    .C(_0293_),
    .Y(_0294_));
 sg13g2_a221oi_1 _0747_ (.B2(_0291_),
    .C1(_0294_),
    .B1(_0281_),
    .A1(_0273_),
    .Y(_0295_),
    .A2(_0278_));
 sg13g2_nand2_1 _0748_ (.Y(_0296_),
    .A(net39),
    .B(_0231_));
 sg13g2_o21ai_1 _0749_ (.B1(_0296_),
    .Y(_0028_),
    .A1(_0231_),
    .A2(_0295_));
 sg13g2_nand2_1 _0750_ (.Y(_0297_),
    .A(net40),
    .B(_0231_));
 sg13g2_o21ai_1 _0751_ (.B1(_0297_),
    .Y(_0029_),
    .A1(_0231_),
    .A2(_0264_));
 sg13g2_mux2_1 _0752_ (.A0(_0239_),
    .A1(net41),
    .S(_0231_),
    .X(_0030_));
 sg13g2_nand2_1 _0753_ (.Y(_0298_),
    .A(net42),
    .B(_0231_));
 sg13g2_o21ai_1 _0754_ (.B1(_0298_),
    .Y(_0031_),
    .A1(_0231_),
    .A2(_0255_));
 sg13g2_buf_4 place259 (.X(net259),
    .A(\genblk1[1].pipe.eps[0][31] ));
 sg13g2_buf_4 place258 (.X(net258),
    .A(\genblk1[2].pipe.eps[0][28] ));
 sg13g2_inv_2 _0757_ (.Y(_0301_),
    .A(net259));
 sg13g2_buf_4 place257 (.X(net257),
    .A(\genblk1[2].pipe.eps[0][29] ));
 sg13g2_buf_4 place256 (.X(net256),
    .A(\genblk1[2].pipe.eps[0][30] ));
 sg13g2_or2_1 _0760_ (.X(_0304_),
    .B(\genblk1[1].pipe.eps[0][29] ),
    .A(net263));
 sg13g2_buf_4 place255 (.X(net255),
    .A(\genblk1[3].pipe.eps[0][28] ));
 sg13g2_tielo _1220__6 (.L_LO(net57));
 sg13g2_nor2_1 _0763_ (.A(net259),
    .B(_0020_),
    .Y(_0307_));
 sg13g2_nor3_1 _0764_ (.A(net261),
    .B(_0304_),
    .C(_0307_),
    .Y(_0308_));
 sg13g2_a21oi_2 _0765_ (.B1(_0308_),
    .Y(_0309_),
    .A2(net261),
    .A1(_0301_));
 sg13g2_nor2_2 _0766_ (.A(\genblk1[1].pipe.eps[0][26] ),
    .B(\genblk1[1].pipe.eps[0][27] ),
    .Y(_0310_));
 sg13g2_or2_1 _0767_ (.X(_0311_),
    .B(_0310_),
    .A(net264));
 sg13g2_buf_4 place254 (.X(net254),
    .A(\genblk1[3].pipe.eps[0][30] ));
 sg13g2_inv_1 _0769_ (.Y(_0313_),
    .A(net262));
 sg13g2_inv_2 _0770_ (.Y(_0314_),
    .A(_0021_));
 sg13g2_inv_1 _0771_ (.Y(_0315_),
    .A(net260));
 sg13g2_nand2_1 _0772_ (.Y(_0316_),
    .A(net263),
    .B(\genblk1[1].pipe.eps[0][29] ));
 sg13g2_o21ai_1 _0773_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0315_),
    .A2(_0304_));
 sg13g2_nand2b_1 _0774_ (.Y(_0318_),
    .B(\genblk1[1].pipe.eps[0][30] ),
    .A_N(_0021_));
 sg13g2_or4_1 _0775_ (.A(net260),
    .B(net263),
    .C(\genblk1[1].pipe.eps[0][29] ),
    .D(_0020_),
    .X(_0319_));
 sg13g2_a21oi_1 _0776_ (.A1(_0318_),
    .A2(_0319_),
    .Y(_0320_),
    .B1(\genblk1[1].pipe.eps[0][31] ));
 sg13g2_a221oi_1 _0777_ (.B2(net259),
    .C1(_0320_),
    .B1(_0317_),
    .A1(_0313_),
    .Y(_0321_),
    .A2(_0314_));
 sg13g2_a21o_1 _0778_ (.A2(_0021_),
    .A1(_0020_),
    .B1(net262),
    .X(_0322_));
 sg13g2_nand3b_1 _0779_ (.B(net263),
    .C(net262),
    .Y(_0323_),
    .A_N(\genblk1[1].pipe.eps[0][31] ));
 sg13g2_o21ai_1 _0780_ (.B1(_0323_),
    .Y(_0324_),
    .A1(net263),
    .A2(_0322_));
 sg13g2_nor2b_1 _0781_ (.A(net261),
    .B_N(_0020_),
    .Y(_0325_));
 sg13g2_o21ai_1 _0782_ (.B1(_0325_),
    .Y(_0326_),
    .A1(net264),
    .A2(_0310_));
 sg13g2_nand2b_1 _0783_ (.Y(_0327_),
    .B(net263),
    .A_N(_0021_));
 sg13g2_a21oi_1 _0784_ (.A1(net260),
    .A2(_0327_),
    .Y(_0328_),
    .B1(net259));
 sg13g2_o21ai_1 _0785_ (.B1(net261),
    .Y(_0329_),
    .A1(net264),
    .A2(net262));
 sg13g2_or3_1 _0786_ (.A(net260),
    .B(net264),
    .C(net262),
    .X(_0330_));
 sg13g2_a21oi_2 _0787_ (.B1(_0301_),
    .Y(_0331_),
    .A2(_0330_),
    .A1(_0329_));
 sg13g2_a221oi_1 _0788_ (.B2(_0328_),
    .C1(_0331_),
    .B1(_0326_),
    .A1(_0315_),
    .Y(_0332_),
    .A2(_0324_));
 sg13g2_o21ai_1 _0789_ (.B1(_0332_),
    .Y(_0333_),
    .A1(_0311_),
    .A2(_0321_));
 sg13g2_buf_4 place253 (.X(net253),
    .A(\genblk1[3].pipe.eps[0][31] ));
 sg13g2_mux2_1 _0791_ (.A0(_0309_),
    .A1(_0310_),
    .S(_0333_),
    .X(_0335_));
 sg13g2_xor2_1 _0792_ (.B(_0335_),
    .A(net264),
    .X(_0336_));
 sg13g2_nor2b_2 _0793_ (.A(\genblk1[1].pipe.eps[0][27] ),
    .B_N(\genblk1[1].pipe.eps[0][26] ),
    .Y(_0337_));
 sg13g2_nor3_1 _0794_ (.A(\genblk1[1].pipe.eps[0][25] ),
    .B(\genblk1[1].pipe.eps[0][24] ),
    .C(\genblk1[1].pipe.eps[0][26] ),
    .Y(_0338_));
 sg13g2_or2_1 _0795_ (.X(_0339_),
    .B(_0338_),
    .A(_0309_));
 sg13g2_mux2_1 _0796_ (.A0(_0022_),
    .A1(\genblk1[1].pipe.eps[0][27] ),
    .S(_0333_),
    .X(_0340_));
 sg13g2_and2_1 _0797_ (.A(_0309_),
    .B(_0338_),
    .X(_0341_));
 sg13g2_a221oi_1 _0798_ (.B2(_0340_),
    .C1(_0341_),
    .B1(_0339_),
    .A1(_0333_),
    .Y(_0342_),
    .A2(_0337_));
 sg13g2_nor2_2 _0799_ (.A(net259),
    .B(net261),
    .Y(_0343_));
 sg13g2_a21oi_1 _0800_ (.A1(_0336_),
    .A2(_0342_),
    .Y(_0344_),
    .B1(_0343_));
 sg13g2_nor2_1 _0801_ (.A(_0336_),
    .B(_0342_),
    .Y(_0345_));
 sg13g2_nand2_1 _0802_ (.Y(_0346_),
    .A(net262),
    .B(_0309_));
 sg13g2_o21ai_1 _0803_ (.B1(_0346_),
    .Y(_0347_),
    .A1(_0314_),
    .A2(_0309_));
 sg13g2_inv_1 _0804_ (.Y(_0348_),
    .A(_0022_));
 sg13g2_nor3_2 _0805_ (.A(net264),
    .B(_0348_),
    .C(_0337_),
    .Y(_0349_));
 sg13g2_xnor2_1 _0806_ (.Y(_0350_),
    .A(_0343_),
    .B(_0349_));
 sg13g2_xnor2_1 _0807_ (.Y(_0351_),
    .A(_0347_),
    .B(_0350_));
 sg13g2_o21ai_1 _0808_ (.B1(_0316_),
    .Y(_0352_),
    .A1(_0021_),
    .A2(_0304_));
 sg13g2_and2_1 _0809_ (.A(_0020_),
    .B(_0343_),
    .X(_0353_));
 sg13g2_nor2_1 _0810_ (.A(_0315_),
    .B(_0327_),
    .Y(_0354_));
 sg13g2_nor3_1 _0811_ (.A(net261),
    .B(net264),
    .C(_0310_),
    .Y(_0355_));
 sg13g2_o21ai_1 _0812_ (.B1(_0301_),
    .Y(_0356_),
    .A1(_0354_),
    .A2(_0355_));
 sg13g2_o21ai_1 _0813_ (.B1(_0356_),
    .Y(_0357_),
    .A1(_0311_),
    .A2(_0321_));
 sg13g2_nor2_1 _0814_ (.A(net260),
    .B(net264),
    .Y(_0358_));
 sg13g2_a22oi_1 _0815_ (.Y(_0359_),
    .B1(_0322_),
    .B2(_0358_),
    .A2(_0314_),
    .A1(net260));
 sg13g2_nor2_1 _0816_ (.A(net263),
    .B(net262),
    .Y(_0360_));
 sg13g2_o21ai_1 _0817_ (.B1(_0360_),
    .Y(_0361_),
    .A1(net261),
    .A2(_0314_));
 sg13g2_mux2_1 _0818_ (.A0(_0359_),
    .A1(_0361_),
    .S(net259),
    .X(_0362_));
 sg13g2_nor2_1 _0819_ (.A(_0349_),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_nor3_1 _0820_ (.A(net259),
    .B(net261),
    .C(_0020_),
    .Y(_0364_));
 sg13g2_nand2_1 _0821_ (.Y(_0365_),
    .A(_0304_),
    .B(_0364_));
 sg13g2_or4_1 _0822_ (.A(_0331_),
    .B(_0349_),
    .C(_0362_),
    .D(_0364_),
    .X(_0366_));
 sg13g2_o21ai_1 _0823_ (.B1(_0366_),
    .Y(_0367_),
    .A1(_0363_),
    .A2(_0365_));
 sg13g2_inv_1 _0824_ (.Y(_0368_),
    .A(_0331_));
 sg13g2_nor2_1 _0825_ (.A(_0368_),
    .B(_0357_),
    .Y(_0369_));
 sg13g2_a221oi_1 _0826_ (.B2(_0367_),
    .C1(_0369_),
    .B1(_0357_),
    .A1(_0352_),
    .Y(_0370_),
    .A2(_0353_));
 sg13g2_and2_1 _0827_ (.A(net259),
    .B(_0317_),
    .X(_0371_));
 sg13g2_nor2_1 _0828_ (.A(net260),
    .B(_0316_),
    .Y(_0372_));
 sg13g2_a21o_1 _0829_ (.A2(_0360_),
    .A1(_0314_),
    .B1(_0372_),
    .X(_0373_));
 sg13g2_or4_1 _0830_ (.A(_0371_),
    .B(_0320_),
    .C(_0333_),
    .D(_0373_),
    .X(_0374_));
 sg13g2_o21ai_1 _0831_ (.B1(_0374_),
    .Y(_0375_),
    .A1(_0351_),
    .A2(_0370_));
 sg13g2_o21ai_1 _0832_ (.B1(_0375_),
    .Y(_0376_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_or2_1 _0833_ (.X(_0377_),
    .B(\genblk1[1].pipe.counter[0] ),
    .A(\genblk1[1].pipe.counter[1] ));
 sg13g2_nor4_2 _0834_ (.A(\genblk1[1].pipe.counter[2] ),
    .B(\genblk1[1].pipe.counter[3] ),
    .C(\genblk1[1].pipe.counter[4] ),
    .Y(_0378_),
    .D(_0377_));
 sg13g2_and2_1 _0835_ (.A(net276),
    .B(\genblk1[1].pipe.state[0] ),
    .X(_0379_));
 sg13g2_buf_4 place263 (.X(net263),
    .A(\genblk1[1].pipe.eps[0][28] ));
 sg13g2_nor2_2 _0837_ (.A(net275),
    .B(_0379_),
    .Y(_0381_));
 sg13g2_nand3_1 _0838_ (.B(_0378_),
    .C(_0381_),
    .A(\genblk1[1].pipe.state[1] ),
    .Y(_0382_));
 sg13g2_buf_4 place252 (.X(net252),
    .A(_0208_));
 sg13g2_mux2_1 _0840_ (.A0(_0376_),
    .A1(net43),
    .S(_0382_),
    .X(_0046_));
 sg13g2_mux2_1 _0841_ (.A0(_0333_),
    .A1(net44),
    .S(_0382_),
    .X(_0047_));
 sg13g2_inv_1 _0842_ (.Y(_0384_),
    .A(_0309_));
 sg13g2_nand2_1 _0843_ (.Y(_0385_),
    .A(net45),
    .B(_0382_));
 sg13g2_o21ai_1 _0844_ (.B1(_0385_),
    .Y(_0048_),
    .A1(_0382_),
    .A2(_0384_));
 sg13g2_nand2_1 _0845_ (.Y(_0386_),
    .A(net46),
    .B(_0382_));
 sg13g2_o21ai_1 _0846_ (.B1(_0386_),
    .Y(_0049_),
    .A1(_0382_),
    .A2(_0343_));
 sg13g2_buf_4 place251 (.X(net251),
    .A(_0214_));
 sg13g2_buf_4 place250 (.X(net250),
    .A(_0218_));
 sg13g2_xor2_1 _0849_ (.B(net257),
    .A(net258),
    .X(_0389_));
 sg13g2_buf_4 place249 (.X(net249),
    .A(_0222_));
 sg13g2_buf_4 place248 (.X(net248),
    .A(_0227_));
 sg13g2_and2_1 _0852_ (.A(\genblk1[2].pipe.eps[0][31] ),
    .B(net256),
    .X(_0392_));
 sg13g2_buf_4 place247 (.X(net247),
    .A(_0379_));
 sg13g2_nor2_1 _0854_ (.A(net258),
    .B(net257),
    .Y(_0394_));
 sg13g2_or2_1 _0855_ (.X(_0395_),
    .B(_0012_),
    .A(\genblk1[2].pipe.eps[0][31] ));
 sg13g2_a21oi_2 _0856_ (.B1(net256),
    .Y(_0396_),
    .A2(_0395_),
    .A1(_0394_));
 sg13g2_nor2_2 _0857_ (.A(_0392_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_mux2_1 _0858_ (.A0(_0389_),
    .A1(_0016_),
    .S(_0397_),
    .X(_0398_));
 sg13g2_inv_1 _0859_ (.Y(_0399_),
    .A(_0016_));
 sg13g2_mux2_1 _0860_ (.A0(\genblk1[2].pipe.eps[0][28] ),
    .A1(\genblk1[2].pipe.eps[0][31] ),
    .S(\genblk1[2].pipe.eps[0][30] ),
    .X(_0400_));
 sg13g2_inv_1 _0861_ (.Y(_0401_),
    .A(net257));
 sg13g2_o21ai_1 _0862_ (.B1(_0401_),
    .Y(_0402_),
    .A1(_0399_),
    .A2(_0400_));
 sg13g2_nor2b_1 _0863_ (.A(_0016_),
    .B_N(net256),
    .Y(_0403_));
 sg13g2_nor3_1 _0864_ (.A(net256),
    .B(net257),
    .C(_0012_),
    .Y(_0404_));
 sg13g2_inv_1 _0865_ (.Y(_0405_),
    .A(\genblk1[2].pipe.eps[0][31] ));
 sg13g2_o21ai_1 _0866_ (.B1(_0405_),
    .Y(_0406_),
    .A1(_0403_),
    .A2(_0404_));
 sg13g2_or2_1 _0867_ (.X(_0407_),
    .B(\genblk1[2].pipe.eps[0][30] ),
    .A(\genblk1[2].pipe.eps[0][31] ));
 sg13g2_buf_4 place246 (.X(net246),
    .A(_0463_));
 sg13g2_inv_2 _0869_ (.Y(_0409_),
    .A(\genblk1[2].pipe.eps[0][28] ));
 sg13g2_nand2b_1 _0870_ (.Y(_0410_),
    .B(_0409_),
    .A_N(_0407_));
 sg13g2_nand3_1 _0871_ (.B(net256),
    .C(net258),
    .A(_0405_),
    .Y(_0411_));
 sg13g2_a22oi_1 _0872_ (.Y(_0412_),
    .B1(_0410_),
    .B2(_0411_),
    .A2(_0406_),
    .A1(_0402_));
 sg13g2_mux2_1 _0873_ (.A0(\genblk1[2].pipe.eps[0][28] ),
    .A1(\genblk1[2].pipe.eps[0][31] ),
    .S(net257),
    .X(_0413_));
 sg13g2_buf_1 output51 (.A(net51),
    .X(valid));
 sg13g2_buf_4 output50 (.X(results[79]),
    .A(net50));
 sg13g2_or3_1 _0876_ (.A(\genblk1[2].pipe.eps[0][26] ),
    .B(\genblk1[2].pipe.eps[0][27] ),
    .C(\genblk1[2].pipe.eps[0][28] ),
    .X(_0416_));
 sg13g2_nor2b_1 _0877_ (.A(_0413_),
    .B_N(_0416_),
    .Y(_0417_));
 sg13g2_nor2_1 _0878_ (.A(\genblk1[2].pipe.eps[0][26] ),
    .B(\genblk1[2].pipe.eps[0][27] ),
    .Y(_0418_));
 sg13g2_a221oi_1 _0879_ (.B2(_0409_),
    .C1(_0413_),
    .B1(_0418_),
    .A1(_0016_),
    .Y(_0419_),
    .A2(_0407_));
 sg13g2_a21o_1 _0880_ (.A2(_0417_),
    .A1(_0392_),
    .B1(_0419_),
    .X(_0420_));
 sg13g2_o21ai_1 _0881_ (.B1(net256),
    .Y(_0421_),
    .A1(net258),
    .A2(net257));
 sg13g2_or3_1 _0882_ (.A(net256),
    .B(net258),
    .C(net257),
    .X(_0422_));
 sg13g2_a21o_2 _0883_ (.A2(_0422_),
    .A1(_0421_),
    .B1(_0405_),
    .X(_0423_));
 sg13g2_o21ai_1 _0884_ (.B1(_0423_),
    .Y(_0424_),
    .A1(_0012_),
    .A2(_0407_));
 sg13g2_nor3_2 _0885_ (.A(_0412_),
    .B(_0420_),
    .C(_0424_),
    .Y(_0425_));
 sg13g2_buf_4 output49 (.X(results[78]),
    .A(net49));
 sg13g2_nand2b_1 _0887_ (.Y(_0427_),
    .B(\genblk1[2].pipe.eps[0][26] ),
    .A_N(\genblk1[2].pipe.eps[0][27] ));
 sg13g2_and3_2 _0888_ (.X(_0428_),
    .A(_0409_),
    .B(_0018_),
    .C(_0427_));
 sg13g2_a21oi_1 _0889_ (.A1(\genblk1[2].pipe.eps[0][31] ),
    .A2(net258),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_nand2_1 _0890_ (.Y(_0430_),
    .A(_0407_),
    .B(_0429_));
 sg13g2_a21o_1 _0891_ (.A2(_0406_),
    .A1(_0402_),
    .B1(_0428_),
    .X(_0431_));
 sg13g2_nand3_1 _0892_ (.B(_0406_),
    .C(_0428_),
    .A(_0402_),
    .Y(_0432_));
 sg13g2_nor2_1 _0893_ (.A(_0012_),
    .B(_0394_),
    .Y(_0433_));
 sg13g2_nor2_1 _0894_ (.A(_0407_),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_nand3_1 _0895_ (.B(_0432_),
    .C(_0434_),
    .A(_0431_),
    .Y(_0435_));
 sg13g2_o21ai_1 _0896_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0398_),
    .A2(_0430_));
 sg13g2_or2_1 _0897_ (.X(_0437_),
    .B(_0420_),
    .A(_0412_));
 sg13g2_or4_1 _0898_ (.A(net256),
    .B(net258),
    .C(net257),
    .D(_0012_),
    .X(_0438_));
 sg13g2_and3_1 _0899_ (.X(_0439_),
    .A(_0437_),
    .B(_0423_),
    .C(_0438_));
 sg13g2_a21oi_1 _0900_ (.A1(_0431_),
    .A2(_0432_),
    .Y(_0440_),
    .B1(_0423_));
 sg13g2_nor2b_1 _0901_ (.A(_0437_),
    .B_N(_0440_),
    .Y(_0441_));
 sg13g2_a221oi_1 _0902_ (.B2(_0439_),
    .C1(_0441_),
    .B1(_0436_),
    .A1(_0398_),
    .Y(_0442_),
    .A2(_0425_));
 sg13g2_nor3_2 _0903_ (.A(\genblk1[2].pipe.eps[0][25] ),
    .B(\genblk1[2].pipe.eps[0][24] ),
    .C(\genblk1[2].pipe.eps[0][26] ),
    .Y(_0443_));
 sg13g2_nand2b_1 _0904_ (.Y(_0444_),
    .B(_0397_),
    .A_N(_0443_));
 sg13g2_mux2_1 _0905_ (.A0(\genblk1[2].pipe.eps[0][27] ),
    .A1(_0018_),
    .S(_0425_),
    .X(_0445_));
 sg13g2_o21ai_1 _0906_ (.B1(\genblk1[2].pipe.eps[0][28] ),
    .Y(_0446_),
    .A1(\genblk1[2].pipe.eps[0][26] ),
    .A2(\genblk1[2].pipe.eps[0][27] ));
 sg13g2_a21o_1 _0907_ (.A2(_0446_),
    .A1(_0416_),
    .B1(_0425_),
    .X(_0447_));
 sg13g2_nor3_1 _0908_ (.A(_0409_),
    .B(_0392_),
    .C(_0396_),
    .Y(_0448_));
 sg13g2_nor2_1 _0909_ (.A(net258),
    .B(_0397_),
    .Y(_0449_));
 sg13g2_o21ai_1 _0910_ (.B1(_0425_),
    .Y(_0450_),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_o21ai_1 _0911_ (.B1(_0443_),
    .Y(_0451_),
    .A1(_0392_),
    .A2(_0396_));
 sg13g2_o21ai_1 _0912_ (.B1(_0451_),
    .Y(_0452_),
    .A1(_0427_),
    .A2(_0425_));
 sg13g2_a221oi_1 _0913_ (.B2(_0450_),
    .C1(_0452_),
    .B1(_0447_),
    .A1(_0444_),
    .Y(_0453_),
    .A2(_0445_));
 sg13g2_a21oi_1 _0914_ (.A1(_0447_),
    .A2(_0450_),
    .Y(_0454_),
    .B1(_0407_));
 sg13g2_inv_1 _0915_ (.Y(_0455_),
    .A(\genblk1[2].pipe.eps[0][27] ));
 sg13g2_nor3_1 _0916_ (.A(_0392_),
    .B(_0396_),
    .C(_0443_),
    .Y(_0456_));
 sg13g2_nor3_1 _0917_ (.A(_0455_),
    .B(_0425_),
    .C(_0456_),
    .Y(_0457_));
 sg13g2_and3_1 _0918_ (.X(_0458_),
    .A(_0018_),
    .B(_0425_),
    .C(_0444_));
 sg13g2_nor4_1 _0919_ (.A(_0407_),
    .B(_0452_),
    .C(_0457_),
    .D(_0458_),
    .Y(_0459_));
 sg13g2_or4_1 _0920_ (.A(_0442_),
    .B(_0453_),
    .C(_0454_),
    .D(_0459_),
    .X(_0460_));
 sg13g2_or2_1 _0921_ (.X(_0461_),
    .B(\genblk1[2].pipe.counter[1] ),
    .A(\genblk1[2].pipe.counter[0] ));
 sg13g2_nor4_2 _0922_ (.A(\genblk1[2].pipe.counter[2] ),
    .B(\genblk1[2].pipe.counter[3] ),
    .C(\genblk1[2].pipe.counter[4] ),
    .Y(_0462_),
    .D(_0461_));
 sg13g2_and2_1 _0923_ (.A(net276),
    .B(\genblk1[2].pipe.state[0] ),
    .X(_0463_));
 sg13g2_buf_2 output48 (.A(net48),
    .X(results[77]));
 sg13g2_nor2_2 _0925_ (.A(net275),
    .B(_0463_),
    .Y(_0465_));
 sg13g2_nand3_1 _0926_ (.B(_0462_),
    .C(_0465_),
    .A(\genblk1[2].pipe.state[1] ),
    .Y(_0466_));
 sg13g2_buf_2 output47 (.A(net47),
    .X(results[76]));
 sg13g2_mux2_1 _0928_ (.A0(_0460_),
    .A1(net47),
    .S(_0466_),
    .X(_0064_));
 sg13g2_nand2_1 _0929_ (.Y(_0468_),
    .A(net48),
    .B(_0466_));
 sg13g2_o21ai_1 _0930_ (.B1(_0468_),
    .Y(_0065_),
    .A1(_0466_),
    .A2(_0425_));
 sg13g2_nand2_1 _0931_ (.Y(_0469_),
    .A(net49),
    .B(_0466_));
 sg13g2_o21ai_1 _0932_ (.B1(_0469_),
    .Y(_0066_),
    .A1(_0466_),
    .A2(_0397_));
 sg13g2_mux2_1 _0933_ (.A0(_0407_),
    .A1(net50),
    .S(_0466_),
    .X(_0067_));
 sg13g2_buf_1 output46 (.A(net46),
    .X(results[47]));
 sg13g2_buf_1 output45 (.A(net45),
    .X(results[46]));
 sg13g2_nor2b_1 _0936_ (.A(net253),
    .B_N(net254),
    .Y(_0472_));
 sg13g2_buf_1 output44 (.A(net44),
    .X(results[45]));
 sg13g2_buf_1 output43 (.A(net43),
    .X(results[44]));
 sg13g2_nor2_1 _0939_ (.A(net253),
    .B(_0015_),
    .Y(_0475_));
 sg13g2_nor4_1 _0940_ (.A(net254),
    .B(net255),
    .C(\genblk1[3].pipe.eps[0][29] ),
    .D(_0475_),
    .Y(_0476_));
 sg13g2_nor2_2 _0941_ (.A(_0472_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nor3_1 _0942_ (.A(\genblk1[3].pipe.eps[0][25] ),
    .B(\genblk1[3].pipe.eps[0][24] ),
    .C(\genblk1[3].pipe.eps[0][26] ),
    .Y(_0478_));
 sg13g2_or2_1 _0943_ (.X(_0479_),
    .B(_0478_),
    .A(_0477_));
 sg13g2_nor2_1 _0944_ (.A(net255),
    .B(\genblk1[3].pipe.eps[0][29] ),
    .Y(_0480_));
 sg13g2_nor2_1 _0945_ (.A(net254),
    .B(_0015_),
    .Y(_0481_));
 sg13g2_nand2_1 _0946_ (.Y(_0482_),
    .A(_0480_),
    .B(_0481_));
 sg13g2_nand2_1 _0947_ (.Y(_0483_),
    .A(\genblk1[3].pipe.eps[0][30] ),
    .B(\genblk1[3].pipe.eps[0][28] ));
 sg13g2_or3_1 _0948_ (.A(net254),
    .B(\genblk1[3].pipe.eps[0][28] ),
    .C(\genblk1[3].pipe.eps[0][29] ),
    .X(_0484_));
 sg13g2_a21o_1 _0949_ (.A2(_0484_),
    .A1(_0483_),
    .B1(_0014_),
    .X(_0485_));
 sg13g2_a21oi_1 _0950_ (.A1(_0482_),
    .A2(_0485_),
    .Y(_0486_),
    .B1(net253));
 sg13g2_nand2b_1 _0951_ (.Y(_0487_),
    .B(_0014_),
    .A_N(\genblk1[3].pipe.eps[0][28] ));
 sg13g2_inv_1 _0952_ (.Y(_0488_),
    .A(\genblk1[3].pipe.eps[0][29] ));
 sg13g2_o21ai_1 _0953_ (.B1(_0488_),
    .Y(_0489_),
    .A1(\genblk1[3].pipe.eps[0][30] ),
    .A2(_0487_));
 sg13g2_nor2_1 _0954_ (.A(\genblk1[3].pipe.eps[0][26] ),
    .B(\genblk1[3].pipe.eps[0][27] ),
    .Y(_0490_));
 sg13g2_mux2_1 _0955_ (.A0(_0490_),
    .A1(_0488_),
    .S(\genblk1[3].pipe.eps[0][28] ),
    .X(_0491_));
 sg13g2_a221oi_1 _0956_ (.B2(_0014_),
    .C1(_0491_),
    .B1(_0472_),
    .A1(net253),
    .Y(_0492_),
    .A2(_0489_));
 sg13g2_o21ai_1 _0957_ (.B1(net254),
    .Y(_0493_),
    .A1(net255),
    .A2(\genblk1[3].pipe.eps[0][29] ));
 sg13g2_inv_1 _0958_ (.Y(_0494_),
    .A(net253));
 sg13g2_a21oi_1 _0959_ (.A1(_0484_),
    .A2(_0493_),
    .Y(_0495_),
    .B1(_0494_));
 sg13g2_nor3_1 _0960_ (.A(net253),
    .B(net254),
    .C(_0015_),
    .Y(_0496_));
 sg13g2_nor4_2 _0961_ (.A(_0486_),
    .B(_0492_),
    .C(_0495_),
    .Y(_0497_),
    .D(_0496_));
 sg13g2_mux2_1 _0962_ (.A0(\genblk1[3].pipe.eps[0][27] ),
    .A1(_0010_),
    .S(_0497_),
    .X(_0498_));
 sg13g2_nand2b_2 _0963_ (.Y(_0499_),
    .B(\genblk1[3].pipe.eps[0][26] ),
    .A_N(\genblk1[3].pipe.eps[0][27] ));
 sg13g2_nand2_1 _0964_ (.Y(_0500_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_o21ai_1 _0965_ (.B1(_0500_),
    .Y(_0501_),
    .A1(_0497_),
    .A2(_0499_));
 sg13g2_a21oi_1 _0966_ (.A1(_0479_),
    .A2(_0498_),
    .Y(_0502_),
    .B1(_0501_));
 sg13g2_mux2_1 _0967_ (.A0(_0490_),
    .A1(_0477_),
    .S(_0497_),
    .X(_0503_));
 sg13g2_xor2_1 _0968_ (.B(_0503_),
    .A(net255),
    .X(_0504_));
 sg13g2_nor2_2 _0969_ (.A(net253),
    .B(net254),
    .Y(_0505_));
 sg13g2_a21oi_1 _0970_ (.A1(_0502_),
    .A2(_0504_),
    .Y(_0506_),
    .B1(_0505_));
 sg13g2_nor2_1 _0971_ (.A(_0502_),
    .B(_0504_),
    .Y(_0507_));
 sg13g2_o21ai_1 _0972_ (.B1(_0505_),
    .Y(_0508_),
    .A1(_0015_),
    .A2(_0480_));
 sg13g2_xor2_1 _0973_ (.B(\genblk1[3].pipe.eps[0][29] ),
    .A(net255),
    .X(_0509_));
 sg13g2_mux2_1 _0974_ (.A0(_0014_),
    .A1(_0509_),
    .S(_0477_),
    .X(_0510_));
 sg13g2_nand2b_1 _0975_ (.Y(_0511_),
    .B(net254),
    .A_N(net253));
 sg13g2_nor2b_1 _0976_ (.A(net255),
    .B_N(_0010_),
    .Y(_0512_));
 sg13g2_a22oi_1 _0977_ (.Y(_0513_),
    .B1(_0499_),
    .B2(_0512_),
    .A2(_0511_),
    .A1(net255));
 sg13g2_xnor2_1 _0978_ (.Y(_0514_),
    .A(_0510_),
    .B(_0513_));
 sg13g2_mux2_1 _0979_ (.A0(_0505_),
    .A1(_0508_),
    .S(_0514_),
    .X(_0515_));
 sg13g2_a21oi_1 _0980_ (.A1(_0480_),
    .A2(_0481_),
    .Y(_0516_),
    .B1(_0495_));
 sg13g2_nor2_1 _0981_ (.A(_0486_),
    .B(_0492_),
    .Y(_0517_));
 sg13g2_nand2b_1 _0982_ (.Y(_0518_),
    .B(_0517_),
    .A_N(_0516_));
 sg13g2_nand2b_1 _0983_ (.Y(_0519_),
    .B(_0513_),
    .A_N(_0505_));
 sg13g2_o21ai_1 _0984_ (.B1(_0519_),
    .Y(_0520_),
    .A1(_0513_),
    .A2(_0508_));
 sg13g2_a221oi_1 _0985_ (.B2(_0512_),
    .C1(_0508_),
    .B1(_0499_),
    .A1(net255),
    .Y(_0521_),
    .A2(_0511_));
 sg13g2_mux2_1 _0986_ (.A0(_0520_),
    .A1(_0521_),
    .S(_0510_),
    .X(_0522_));
 sg13g2_nor2b_1 _0987_ (.A(_0517_),
    .B_N(_0516_),
    .Y(_0523_));
 sg13g2_a22oi_1 _0988_ (.Y(_0524_),
    .B1(_0522_),
    .B2(_0523_),
    .A2(_0510_),
    .A1(_0497_));
 sg13g2_o21ai_1 _0989_ (.B1(_0524_),
    .Y(_0525_),
    .A1(_0515_),
    .A2(_0518_));
 sg13g2_o21ai_1 _0990_ (.B1(_0525_),
    .Y(_0526_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_inv_1 _0991_ (.Y(_0527_),
    .A(net271));
 sg13g2_inv_1 _0992_ (.Y(_0528_),
    .A(\genblk1[3].pipe.counter[4] ));
 sg13g2_or2_1 _0993_ (.X(_0529_),
    .B(\genblk1[3].pipe.counter[1] ),
    .A(\genblk1[3].pipe.counter[0] ));
 sg13g2_nor2_1 _0994_ (.A(\genblk1[3].pipe.counter[2] ),
    .B(_0529_),
    .Y(_0530_));
 sg13g2_nand2_1 _0995_ (.Y(_0531_),
    .A(\genblk1[3].pipe.state[1] ),
    .B(_0530_));
 sg13g2_nor2_1 _0996_ (.A(\genblk1[3].pipe.counter[3] ),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nand4_1 _0997_ (.B(_0528_),
    .C(_0222_),
    .A(_0527_),
    .Y(_0533_),
    .D(_0532_));
 sg13g2_buf_1 output42 (.A(net42),
    .X(results[15]));
 sg13g2_mux2_1 _0999_ (.A0(_0526_),
    .A1(net35),
    .S(_0533_),
    .X(_0082_));
 sg13g2_nand2_1 _1000_ (.Y(_0535_),
    .A(net36),
    .B(_0533_));
 sg13g2_o21ai_1 _1001_ (.B1(_0535_),
    .Y(_0083_),
    .A1(_0533_),
    .A2(_0497_));
 sg13g2_mux2_1 _1002_ (.A0(_0477_),
    .A1(net37),
    .S(_0533_),
    .X(_0084_));
 sg13g2_nand2_1 _1003_ (.Y(_0536_),
    .A(net38),
    .B(_0533_));
 sg13g2_o21ai_1 _1004_ (.B1(_0536_),
    .Y(_0085_),
    .A1(_0533_),
    .A2(_0505_));
 sg13g2_nor3_1 _1005_ (.A(\genblk1[0].pipe.counter[1] ),
    .B(\genblk1[0].pipe.counter[0] ),
    .C(\genblk1[0].pipe.counter[2] ),
    .Y(_0537_));
 sg13g2_a21o_1 _1006_ (.A2(_0537_),
    .A1(_0230_),
    .B1(_0213_),
    .X(_0538_));
 sg13g2_buf_2 output41 (.A(net41),
    .X(results[14]));
 sg13g2_or2_1 _1008_ (.X(_0540_),
    .B(_0538_),
    .A(\genblk1[0].pipe.counter[0] ));
 sg13g2_a21oi_1 _1009_ (.A1(_0213_),
    .A2(\genblk1[0].pipe.counter[0] ),
    .Y(_0541_),
    .B1(_0227_));
 sg13g2_a21oi_1 _1010_ (.A1(_0540_),
    .A2(_0541_),
    .Y(_0023_),
    .B1(net34));
 sg13g2_xor2_1 _1011_ (.B(_0540_),
    .A(\genblk1[0].pipe.counter[1] ),
    .X(_0542_));
 sg13g2_a21oi_1 _1012_ (.A1(_0214_),
    .A2(_0542_),
    .Y(_0024_),
    .B1(net34));
 sg13g2_nor2_1 _1013_ (.A(\genblk1[0].pipe.counter[2] ),
    .B(_0230_),
    .Y(_0543_));
 sg13g2_mux2_1 _1014_ (.A0(\genblk1[0].pipe.counter[2] ),
    .A1(_0543_),
    .S(_0225_),
    .X(_0544_));
 sg13g2_and2_1 _1015_ (.A(_0229_),
    .B(_0544_),
    .X(_0025_));
 sg13g2_nor2b_1 _1016_ (.A(\genblk1[0].pipe.counter[3] ),
    .B_N(\genblk1[0].pipe.counter[4] ),
    .Y(_0545_));
 sg13g2_mux2_1 _1017_ (.A0(\genblk1[0].pipe.counter[3] ),
    .A1(_0545_),
    .S(_0226_),
    .X(_0546_));
 sg13g2_and2_1 _1018_ (.A(_0229_),
    .B(_0546_),
    .X(_0026_));
 sg13g2_nand2b_1 _1019_ (.Y(_0547_),
    .B(_0226_),
    .A_N(\genblk1[0].pipe.counter[3] ));
 sg13g2_and3_1 _1020_ (.X(_0027_),
    .A(\genblk1[0].pipe.counter[4] ),
    .B(_0229_),
    .C(_0547_));
 sg13g2_buf_1 output40 (.A(net40),
    .X(results[13]));
 sg13g2_buf_4 output39 (.X(results[12]),
    .A(net39));
 sg13g2_buf_4 output38 (.X(results[111]),
    .A(net38));
 sg13g2_buf_8 output37 (.A(net37),
    .X(results[110]));
 sg13g2_buf_4 output36 (.X(results[109]),
    .A(net36));
 sg13g2_buf_4 output35 (.X(results[108]),
    .A(net35));
 sg13g2_nand2_1 _1027_ (.Y(_0554_),
    .A(net9),
    .B(net248));
 sg13g2_nand3_1 _1028_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][24] ),
    .Y(_0555_));
 sg13g2_a21oi_1 _1029_ (.A1(_0554_),
    .A2(_0555_),
    .Y(_0032_),
    .B1(net268));
 sg13g2_nand2_1 _1030_ (.Y(_0556_),
    .A(net10),
    .B(net248));
 sg13g2_nand3_1 _1031_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][25] ),
    .Y(_0557_));
 sg13g2_a21oi_1 _1032_ (.A1(_0556_),
    .A2(_0557_),
    .Y(_0033_),
    .B1(net268));
 sg13g2_nand2_1 _1033_ (.Y(_0558_),
    .A(net11),
    .B(net248));
 sg13g2_nand3_1 _1034_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][26] ),
    .Y(_0559_));
 sg13g2_a21oi_1 _1035_ (.A1(_0558_),
    .A2(_0559_),
    .Y(_0034_),
    .B1(net268));
 sg13g2_nand2_1 _1036_ (.Y(_0560_),
    .A(net12),
    .B(net248));
 sg13g2_nand3_1 _1037_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][27] ),
    .Y(_0561_));
 sg13g2_a21oi_1 _1038_ (.A1(_0560_),
    .A2(_0561_),
    .Y(_0035_),
    .B1(net268));
 sg13g2_nand2_1 _1039_ (.Y(_0562_),
    .A(net13),
    .B(net248));
 sg13g2_buf_8 input34 (.A(reset),
    .X(net34));
 sg13g2_nand3_1 _1041_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][28] ),
    .Y(_0564_));
 sg13g2_a21oi_1 _1042_ (.A1(_0562_),
    .A2(_0564_),
    .Y(_0036_),
    .B1(net268));
 sg13g2_nand2_1 _1043_ (.Y(_0565_),
    .A(net14),
    .B(net248));
 sg13g2_nand3_1 _1044_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][29] ),
    .Y(_0566_));
 sg13g2_a21oi_1 _1045_ (.A1(_0565_),
    .A2(_0566_),
    .Y(_0037_),
    .B1(net268));
 sg13g2_buf_1 input33 (.A(ready),
    .X(net33));
 sg13g2_nand2_1 _1047_ (.Y(_0568_),
    .A(net15),
    .B(net248));
 sg13g2_nand3_1 _1048_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][30] ),
    .Y(_0569_));
 sg13g2_buf_1 input32 (.A(queries[95]),
    .X(net32));
 sg13g2_a21oi_1 _1050_ (.A1(_0568_),
    .A2(_0569_),
    .Y(_0038_),
    .B1(net268));
 sg13g2_nand2_1 _1051_ (.Y(_0571_),
    .A(net16),
    .B(net248));
 sg13g2_nand3_1 _1052_ (.B(net251),
    .C(net244),
    .A(\genblk1[0].pipe.eps[0][31] ),
    .Y(_0572_));
 sg13g2_a21oi_1 _1053_ (.A1(_0571_),
    .A2(_0572_),
    .Y(_0039_),
    .B1(net268));
 sg13g2_inv_1 _1054_ (.Y(_0573_),
    .A(\genblk1[0].pipe.valid ));
 sg13g2_o21ai_1 _1055_ (.B1(_0231_),
    .Y(_0040_),
    .A1(_0573_),
    .A2(net273));
 sg13g2_or2_1 _1056_ (.X(_0574_),
    .B(_0378_),
    .A(_0019_));
 sg13g2_buf_1 input31 (.A(queries[94]),
    .X(net31));
 sg13g2_or2_1 _1058_ (.X(_0576_),
    .B(_0574_),
    .A(\genblk1[1].pipe.counter[0] ));
 sg13g2_a21oi_1 _1059_ (.A1(\genblk1[1].pipe.counter[0] ),
    .A2(_0019_),
    .Y(_0577_),
    .B1(_0379_));
 sg13g2_a21oi_1 _1060_ (.A1(_0576_),
    .A2(_0577_),
    .Y(_0041_),
    .B1(net275));
 sg13g2_xor2_1 _1061_ (.B(_0576_),
    .A(\genblk1[1].pipe.counter[1] ),
    .X(_0578_));
 sg13g2_buf_1 input30 (.A(queries[93]),
    .X(net30));
 sg13g2_a21oi_1 _1063_ (.A1(_0218_),
    .A2(_0578_),
    .Y(_0042_),
    .B1(net275));
 sg13g2_nor2_1 _1064_ (.A(_0377_),
    .B(_0574_),
    .Y(_0095_));
 sg13g2_xor2_1 _1065_ (.B(_0095_),
    .A(\genblk1[1].pipe.counter[2] ),
    .X(_0096_));
 sg13g2_and2_1 _1066_ (.A(_0381_),
    .B(_0096_),
    .X(_0043_));
 sg13g2_nor2b_1 _1067_ (.A(\genblk1[1].pipe.counter[3] ),
    .B_N(\genblk1[1].pipe.counter[4] ),
    .Y(_0097_));
 sg13g2_nor3_1 _1068_ (.A(\genblk1[1].pipe.counter[2] ),
    .B(_0019_),
    .C(_0377_),
    .Y(_0098_));
 sg13g2_mux2_1 _1069_ (.A0(\genblk1[1].pipe.counter[3] ),
    .A1(_0097_),
    .S(_0098_),
    .X(_0099_));
 sg13g2_and2_1 _1070_ (.A(_0381_),
    .B(_0099_),
    .X(_0044_));
 sg13g2_nand2b_1 _1071_ (.Y(_0100_),
    .B(_0098_),
    .A_N(\genblk1[1].pipe.counter[3] ));
 sg13g2_and3_1 _1072_ (.X(_0045_),
    .A(\genblk1[1].pipe.counter[4] ),
    .B(_0381_),
    .C(_0100_));
 sg13g2_buf_1 input29 (.A(queries[92]),
    .X(net29));
 sg13g2_buf_1 input28 (.A(queries[91]),
    .X(net28));
 sg13g2_buf_1 input27 (.A(queries[90]),
    .X(net27));
 sg13g2_buf_1 input26 (.A(queries[89]),
    .X(net26));
 sg13g2_buf_1 input25 (.A(queries[88]),
    .X(net25));
 sg13g2_nand2_1 _1078_ (.Y(_0106_),
    .A(net17),
    .B(net247));
 sg13g2_nand3_1 _1079_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][24] ),
    .Y(_0107_));
 sg13g2_a21oi_1 _1080_ (.A1(_0106_),
    .A2(_0107_),
    .Y(_0050_),
    .B1(net272));
 sg13g2_nand2_1 _1081_ (.Y(_0108_),
    .A(net18),
    .B(net247));
 sg13g2_nand3_1 _1082_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][25] ),
    .Y(_0109_));
 sg13g2_a21oi_1 _1083_ (.A1(_0108_),
    .A2(_0109_),
    .Y(_0051_),
    .B1(net272));
 sg13g2_nand2_1 _1084_ (.Y(_0110_),
    .A(net19),
    .B(net247));
 sg13g2_nand3_1 _1085_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][26] ),
    .Y(_0111_));
 sg13g2_a21oi_1 _1086_ (.A1(_0110_),
    .A2(_0111_),
    .Y(_0052_),
    .B1(net272));
 sg13g2_nand2_1 _1087_ (.Y(_0112_),
    .A(net20),
    .B(net247));
 sg13g2_buf_1 input24 (.A(queries[63]),
    .X(net24));
 sg13g2_nand3_1 _1089_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][27] ),
    .Y(_0114_));
 sg13g2_a21oi_1 _1090_ (.A1(_0112_),
    .A2(_0114_),
    .Y(_0053_),
    .B1(net272));
 sg13g2_nand2_1 _1091_ (.Y(_0115_),
    .A(net21),
    .B(net247));
 sg13g2_nand3_1 _1092_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][28] ),
    .Y(_0116_));
 sg13g2_a21oi_1 _1093_ (.A1(_0115_),
    .A2(_0116_),
    .Y(_0054_),
    .B1(net272));
 sg13g2_nand2_1 _1094_ (.Y(_0117_),
    .A(net22),
    .B(net247));
 sg13g2_nand3_1 _1095_ (.B(net250),
    .C(net243),
    .A(net262),
    .Y(_0118_));
 sg13g2_buf_1 input23 (.A(queries[62]),
    .X(net23));
 sg13g2_a21oi_1 _1097_ (.A1(_0117_),
    .A2(_0118_),
    .Y(_0055_),
    .B1(net272));
 sg13g2_buf_1 input22 (.A(queries[61]),
    .X(net22));
 sg13g2_nand2_1 _1099_ (.Y(_0121_),
    .A(net23),
    .B(net247));
 sg13g2_nand3_1 _1100_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][30] ),
    .Y(_0122_));
 sg13g2_a21oi_1 _1101_ (.A1(_0121_),
    .A2(_0122_),
    .Y(_0056_),
    .B1(net272));
 sg13g2_nand2_1 _1102_ (.Y(_0123_),
    .A(net24),
    .B(net247));
 sg13g2_nand3_1 _1103_ (.B(net250),
    .C(net243),
    .A(\genblk1[1].pipe.eps[0][31] ),
    .Y(_0124_));
 sg13g2_a21oi_1 _1104_ (.A1(_0123_),
    .A2(_0124_),
    .Y(_0057_),
    .B1(net272));
 sg13g2_buf_1 input21 (.A(queries[60]),
    .X(net21));
 sg13g2_nor2_1 _1106_ (.A(_0019_),
    .B(_0379_),
    .Y(_0126_));
 sg13g2_a21oi_1 _1107_ (.A1(_0378_),
    .A2(_0126_),
    .Y(_0127_),
    .B1(\genblk1[1].pipe.valid ));
 sg13g2_nor2_1 _1108_ (.A(net275),
    .B(_0127_),
    .Y(_0058_));
 sg13g2_or2_1 _1109_ (.X(_0128_),
    .B(_0462_),
    .A(_0009_));
 sg13g2_buf_1 input20 (.A(queries[59]),
    .X(net20));
 sg13g2_or2_1 _1111_ (.X(_0130_),
    .B(_0128_),
    .A(\genblk1[2].pipe.counter[0] ));
 sg13g2_a21oi_1 _1112_ (.A1(\genblk1[2].pipe.counter[0] ),
    .A2(_0009_),
    .Y(_0131_),
    .B1(_0463_));
 sg13g2_a21oi_1 _1113_ (.A1(_0130_),
    .A2(_0131_),
    .Y(_0059_),
    .B1(net273));
 sg13g2_xor2_1 _1114_ (.B(_0130_),
    .A(\genblk1[2].pipe.counter[1] ),
    .X(_0132_));
 sg13g2_a21oi_1 _1115_ (.A1(_0208_),
    .A2(_0132_),
    .Y(_0060_),
    .B1(net273));
 sg13g2_nor2_1 _1116_ (.A(_0461_),
    .B(_0128_),
    .Y(_0133_));
 sg13g2_xor2_1 _1117_ (.B(_0133_),
    .A(\genblk1[2].pipe.counter[2] ),
    .X(_0134_));
 sg13g2_and2_1 _1118_ (.A(_0465_),
    .B(_0134_),
    .X(_0061_));
 sg13g2_nor2b_1 _1119_ (.A(\genblk1[2].pipe.counter[3] ),
    .B_N(\genblk1[2].pipe.counter[4] ),
    .Y(_0135_));
 sg13g2_nor3_1 _1120_ (.A(\genblk1[2].pipe.counter[2] ),
    .B(_0009_),
    .C(_0461_),
    .Y(_0136_));
 sg13g2_mux2_1 _1121_ (.A0(\genblk1[2].pipe.counter[3] ),
    .A1(_0135_),
    .S(_0136_),
    .X(_0137_));
 sg13g2_and2_1 _1122_ (.A(_0465_),
    .B(_0137_),
    .X(_0062_));
 sg13g2_nand2b_1 _1123_ (.Y(_0138_),
    .B(_0136_),
    .A_N(\genblk1[2].pipe.counter[3] ));
 sg13g2_and3_1 _1124_ (.X(_0063_),
    .A(\genblk1[2].pipe.counter[4] ),
    .B(_0465_),
    .C(_0138_));
 sg13g2_buf_1 input19 (.A(queries[58]),
    .X(net19));
 sg13g2_buf_1 input18 (.A(queries[57]),
    .X(net18));
 sg13g2_buf_1 input17 (.A(queries[56]),
    .X(net17));
 sg13g2_buf_1 input16 (.A(queries[31]),
    .X(net16));
 sg13g2_buf_1 input15 (.A(queries[30]),
    .X(net15));
 sg13g2_nand2_1 _1130_ (.Y(_0144_),
    .A(net25),
    .B(net246));
 sg13g2_nand3_1 _1131_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][24] ),
    .Y(_0145_));
 sg13g2_a21oi_1 _1132_ (.A1(_0144_),
    .A2(_0145_),
    .Y(_0068_),
    .B1(net274));
 sg13g2_nand2_1 _1133_ (.Y(_0146_),
    .A(net26),
    .B(net246));
 sg13g2_nand3_1 _1134_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][25] ),
    .Y(_0147_));
 sg13g2_a21oi_1 _1135_ (.A1(_0146_),
    .A2(_0147_),
    .Y(_0069_),
    .B1(net274));
 sg13g2_nand2_1 _1136_ (.Y(_0148_),
    .A(net27),
    .B(net246));
 sg13g2_nand3_1 _1137_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][26] ),
    .Y(_0149_));
 sg13g2_buf_1 input14 (.A(queries[29]),
    .X(net14));
 sg13g2_a21oi_1 _1139_ (.A1(_0148_),
    .A2(_0149_),
    .Y(_0070_),
    .B1(net274));
 sg13g2_nand2_1 _1140_ (.Y(_0151_),
    .A(net28),
    .B(net246));
 sg13g2_buf_1 input13 (.A(queries[28]),
    .X(net13));
 sg13g2_nand3_1 _1142_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][27] ),
    .Y(_0153_));
 sg13g2_a21oi_1 _1143_ (.A1(_0151_),
    .A2(_0153_),
    .Y(_0071_),
    .B1(net274));
 sg13g2_nand2_1 _1144_ (.Y(_0154_),
    .A(net29),
    .B(net246));
 sg13g2_nand3_1 _1145_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][28] ),
    .Y(_0155_));
 sg13g2_a21oi_1 _1146_ (.A1(_0154_),
    .A2(_0155_),
    .Y(_0072_),
    .B1(net274));
 sg13g2_nand2_1 _1147_ (.Y(_0156_),
    .A(net30),
    .B(net246));
 sg13g2_nand3_1 _1148_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][29] ),
    .Y(_0157_));
 sg13g2_a21oi_1 _1149_ (.A1(_0156_),
    .A2(_0157_),
    .Y(_0073_),
    .B1(net274));
 sg13g2_buf_1 input12 (.A(queries[27]),
    .X(net12));
 sg13g2_nand2_1 _1151_ (.Y(_0159_),
    .A(net31),
    .B(net246));
 sg13g2_nand3_1 _1152_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][30] ),
    .Y(_0160_));
 sg13g2_a21oi_1 _1153_ (.A1(_0159_),
    .A2(_0160_),
    .Y(_0074_),
    .B1(net274));
 sg13g2_nand2_1 _1154_ (.Y(_0161_),
    .A(net32),
    .B(net246));
 sg13g2_nand3_1 _1155_ (.B(net252),
    .C(net242),
    .A(\genblk1[2].pipe.eps[0][31] ),
    .Y(_0162_));
 sg13g2_a21oi_1 _1156_ (.A1(_0161_),
    .A2(_0162_),
    .Y(_0075_),
    .B1(net274));
 sg13g2_buf_1 input11 (.A(queries[26]),
    .X(net11));
 sg13g2_nor2_1 _1158_ (.A(_0009_),
    .B(_0463_),
    .Y(_0164_));
 sg13g2_a21oi_1 _1159_ (.A1(_0462_),
    .A2(_0164_),
    .Y(_0165_),
    .B1(\genblk1[2].pipe.valid ));
 sg13g2_nor2_1 _1160_ (.A(net273),
    .B(_0165_),
    .Y(_0076_));
 sg13g2_nor2_1 _1161_ (.A(\genblk1[3].pipe.counter[3] ),
    .B(\genblk1[3].pipe.counter[4] ),
    .Y(_0166_));
 sg13g2_a21o_2 _1162_ (.A2(_0166_),
    .A1(_0530_),
    .B1(_0221_),
    .X(_0167_));
 sg13g2_buf_1 input10 (.A(queries[25]),
    .X(net10));
 sg13g2_or2_1 _1164_ (.X(_0169_),
    .B(_0167_),
    .A(\genblk1[3].pipe.counter[0] ));
 sg13g2_and2_1 _1165_ (.A(\genblk1[3].pipe.state[0] ),
    .B(net276),
    .X(_0170_));
 sg13g2_buf_1 input9 (.A(queries[24]),
    .X(net9));
 sg13g2_a21oi_1 _1167_ (.A1(_0221_),
    .A2(\genblk1[3].pipe.counter[0] ),
    .Y(_0172_),
    .B1(_0170_));
 sg13g2_a21oi_1 _1168_ (.A1(_0169_),
    .A2(_0172_),
    .Y(_0077_),
    .B1(net271));
 sg13g2_xor2_1 _1169_ (.B(_0169_),
    .A(\genblk1[3].pipe.counter[1] ),
    .X(_0173_));
 sg13g2_a21oi_1 _1170_ (.A1(_0222_),
    .A2(_0173_),
    .Y(_0078_),
    .B1(net271));
 sg13g2_nand2_1 _1171_ (.Y(_0174_),
    .A(_0527_),
    .B(_0222_));
 sg13g2_nor2_1 _1172_ (.A(_0529_),
    .B(_0167_),
    .Y(_0175_));
 sg13g2_xnor2_1 _1173_ (.Y(_0176_),
    .A(\genblk1[3].pipe.counter[2] ),
    .B(_0175_));
 sg13g2_nor2_1 _1174_ (.A(_0174_),
    .B(_0176_),
    .Y(_0079_));
 sg13g2_nor3_1 _1175_ (.A(\genblk1[3].pipe.counter[3] ),
    .B(_0528_),
    .C(_0531_),
    .Y(_0177_));
 sg13g2_a21oi_1 _1176_ (.A1(\genblk1[3].pipe.counter[3] ),
    .A2(_0531_),
    .Y(_0178_),
    .B1(_0177_));
 sg13g2_nor2_1 _1177_ (.A(_0174_),
    .B(_0178_),
    .Y(_0080_));
 sg13g2_nor3_1 _1178_ (.A(_0528_),
    .B(_0532_),
    .C(_0174_),
    .Y(_0081_));
 sg13g2_buf_1 input8 (.A(queries[127]),
    .X(net8));
 sg13g2_buf_1 input7 (.A(queries[126]),
    .X(net7));
 sg13g2_buf_1 input6 (.A(queries[125]),
    .X(net6));
 sg13g2_buf_1 input5 (.A(queries[124]),
    .X(net5));
 sg13g2_nand2_1 _1183_ (.Y(_0183_),
    .A(net1),
    .B(net245));
 sg13g2_nand3_1 _1184_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][24] ),
    .Y(_0184_));
 sg13g2_buf_1 input4 (.A(queries[123]),
    .X(net4));
 sg13g2_a21oi_1 _1186_ (.A1(_0183_),
    .A2(_0184_),
    .Y(_0086_),
    .B1(net269));
 sg13g2_nand2_1 _1187_ (.Y(_0186_),
    .A(net2),
    .B(net245));
 sg13g2_nand3_1 _1188_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][25] ),
    .Y(_0187_));
 sg13g2_a21oi_1 _1189_ (.A1(_0186_),
    .A2(_0187_),
    .Y(_0087_),
    .B1(net269));
 sg13g2_nand2_1 _1190_ (.Y(_0188_),
    .A(net3),
    .B(net245));
 sg13g2_nand3_1 _1191_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][26] ),
    .Y(_0189_));
 sg13g2_a21oi_1 _1192_ (.A1(_0188_),
    .A2(_0189_),
    .Y(_0088_),
    .B1(net269));
 sg13g2_nand2_1 _1193_ (.Y(_0190_),
    .A(net4),
    .B(net245));
 sg13g2_buf_1 input3 (.A(queries[122]),
    .X(net3));
 sg13g2_nand3_1 _1195_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][27] ),
    .Y(_0192_));
 sg13g2_a21oi_1 _1196_ (.A1(_0190_),
    .A2(_0192_),
    .Y(_0089_),
    .B1(net269));
 sg13g2_nand2_1 _1197_ (.Y(_0193_),
    .A(net5),
    .B(net245));
 sg13g2_nand3_1 _1198_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][28] ),
    .Y(_0194_));
 sg13g2_a21oi_1 _1199_ (.A1(_0193_),
    .A2(_0194_),
    .Y(_0090_),
    .B1(net269));
 sg13g2_nand2_1 _1200_ (.Y(_0195_),
    .A(net6),
    .B(net245));
 sg13g2_nand3_1 _1201_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][29] ),
    .Y(_0196_));
 sg13g2_a21oi_1 _1202_ (.A1(_0195_),
    .A2(_0196_),
    .Y(_0091_),
    .B1(net269));
 sg13g2_buf_1 input2 (.A(queries[121]),
    .X(net2));
 sg13g2_nand2_1 _1204_ (.Y(_0198_),
    .A(net7),
    .B(net245));
 sg13g2_nand3_1 _1205_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][30] ),
    .Y(_0199_));
 sg13g2_a21oi_1 _1206_ (.A1(_0198_),
    .A2(_0199_),
    .Y(_0092_),
    .B1(net269));
 sg13g2_nand2_1 _1207_ (.Y(_0200_),
    .A(net8),
    .B(net245));
 sg13g2_nand3_1 _1208_ (.B(net249),
    .C(net241),
    .A(\genblk1[3].pipe.eps[0][31] ),
    .Y(_0201_));
 sg13g2_a21oi_1 _1209_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0093_),
    .B1(net269));
 sg13g2_inv_1 _1210_ (.Y(_0202_),
    .A(\genblk1[3].pipe.valid ));
 sg13g2_o21ai_1 _1211_ (.B1(_0533_),
    .Y(_0094_),
    .A1(_0202_),
    .A2(net271));
 sg13g2_or4_1 _1212_ (.A(\genblk1[1].pipe.valid ),
    .B(\genblk1[0].pipe.valid ),
    .C(\genblk1[3].pipe.valid ),
    .D(\genblk1[2].pipe.valid ),
    .X(net51));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \genblk1[0].pipe.counter[0]$_SDFFE_PP0P__113  (.L_HI(net164));
 sg13g2_buf_1 input1 (.A(queries[120]),
    .X(net1));
 sg13g2_buf_1 _1216_ (.A(net53),
    .X(results[1]));
 sg13g2_buf_1 _1217_ (.A(net54),
    .X(results[2]));
 sg13g2_buf_1 _1218_ (.A(net55),
    .X(results[3]));
 sg13g2_buf_1 _1219_ (.A(net56),
    .X(results[4]));
 sg13g2_buf_1 _1220_ (.A(net57),
    .X(results[5]));
 sg13g2_buf_1 _1221_ (.A(net58),
    .X(results[6]));
 sg13g2_buf_1 _1222_ (.A(net59),
    .X(results[7]));
 sg13g2_buf_1 _1223_ (.A(net60),
    .X(results[8]));
 sg13g2_buf_1 _1224_ (.A(net61),
    .X(results[9]));
 sg13g2_buf_1 _1225_ (.A(net62),
    .X(results[10]));
 sg13g2_buf_1 _1226_ (.A(net63),
    .X(results[11]));
 sg13g2_buf_1 _1227_ (.A(net64),
    .X(results[16]));
 sg13g2_buf_1 _1228_ (.A(net65),
    .X(results[17]));
 sg13g2_buf_1 _1229_ (.A(net66),
    .X(results[18]));
 sg13g2_buf_1 _1230_ (.A(net67),
    .X(results[19]));
 sg13g2_buf_1 _1231_ (.A(net68),
    .X(results[20]));
 sg13g2_buf_1 _1232_ (.A(net69),
    .X(results[21]));
 sg13g2_buf_1 _1233_ (.A(net70),
    .X(results[22]));
 sg13g2_buf_1 _1234_ (.A(net71),
    .X(results[23]));
 sg13g2_buf_1 _1235_ (.A(net72),
    .X(results[24]));
 sg13g2_buf_1 _1236_ (.A(net73),
    .X(results[25]));
 sg13g2_buf_1 _1237_ (.A(net74),
    .X(results[26]));
 sg13g2_buf_1 _1238_ (.A(net75),
    .X(results[27]));
 sg13g2_buf_1 _1239_ (.A(net76),
    .X(results[28]));
 sg13g2_buf_1 _1240_ (.A(net77),
    .X(results[29]));
 sg13g2_buf_1 _1241_ (.A(net78),
    .X(results[30]));
 sg13g2_buf_1 _1242_ (.A(net79),
    .X(results[31]));
 sg13g2_buf_1 _1243_ (.A(net80),
    .X(results[32]));
 sg13g2_buf_1 _1244_ (.A(net81),
    .X(results[33]));
 sg13g2_buf_1 _1245_ (.A(net82),
    .X(results[34]));
 sg13g2_buf_1 _1246_ (.A(net83),
    .X(results[35]));
 sg13g2_buf_1 _1247_ (.A(net84),
    .X(results[36]));
 sg13g2_buf_1 _1248_ (.A(net85),
    .X(results[37]));
 sg13g2_buf_1 _1249_ (.A(net86),
    .X(results[38]));
 sg13g2_buf_1 _1250_ (.A(net87),
    .X(results[39]));
 sg13g2_buf_1 _1251_ (.A(net88),
    .X(results[40]));
 sg13g2_buf_1 _1252_ (.A(net89),
    .X(results[41]));
 sg13g2_buf_1 _1253_ (.A(net90),
    .X(results[42]));
 sg13g2_buf_1 _1254_ (.A(net91),
    .X(results[43]));
 sg13g2_buf_1 _1255_ (.A(net92),
    .X(results[48]));
 sg13g2_buf_1 _1256_ (.A(net93),
    .X(results[49]));
 sg13g2_buf_1 _1257_ (.A(net94),
    .X(results[50]));
 sg13g2_buf_1 _1258_ (.A(net95),
    .X(results[51]));
 sg13g2_buf_1 _1259_ (.A(net96),
    .X(results[52]));
 sg13g2_buf_1 _1260_ (.A(net97),
    .X(results[53]));
 sg13g2_buf_1 _1261_ (.A(net98),
    .X(results[54]));
 sg13g2_buf_1 _1262_ (.A(net99),
    .X(results[55]));
 sg13g2_buf_1 _1263_ (.A(net100),
    .X(results[56]));
 sg13g2_buf_1 _1264_ (.A(net101),
    .X(results[57]));
 sg13g2_buf_1 _1265_ (.A(net102),
    .X(results[58]));
 sg13g2_buf_1 _1266_ (.A(net103),
    .X(results[59]));
 sg13g2_buf_1 _1267_ (.A(net104),
    .X(results[60]));
 sg13g2_buf_1 _1268_ (.A(net105),
    .X(results[61]));
 sg13g2_buf_1 _1269_ (.A(net106),
    .X(results[62]));
 sg13g2_buf_1 _1270_ (.A(net107),
    .X(results[63]));
 sg13g2_buf_1 _1271_ (.A(net108),
    .X(results[64]));
 sg13g2_buf_1 _1272_ (.A(net109),
    .X(results[65]));
 sg13g2_buf_1 _1273_ (.A(net110),
    .X(results[66]));
 sg13g2_buf_1 _1274_ (.A(net111),
    .X(results[67]));
 sg13g2_buf_1 _1275_ (.A(net112),
    .X(results[68]));
 sg13g2_buf_1 _1276_ (.A(net113),
    .X(results[69]));
 sg13g2_buf_1 _1277_ (.A(net114),
    .X(results[70]));
 sg13g2_buf_1 _1278_ (.A(net115),
    .X(results[71]));
 sg13g2_buf_1 _1279_ (.A(net116),
    .X(results[72]));
 sg13g2_buf_1 _1280_ (.A(net117),
    .X(results[73]));
 sg13g2_buf_1 _1281_ (.A(net118),
    .X(results[74]));
 sg13g2_buf_1 _1282_ (.A(net119),
    .X(results[75]));
 sg13g2_buf_1 _1283_ (.A(net120),
    .X(results[80]));
 sg13g2_buf_1 _1284_ (.A(net121),
    .X(results[81]));
 sg13g2_buf_1 _1285_ (.A(net122),
    .X(results[82]));
 sg13g2_buf_1 _1286_ (.A(net123),
    .X(results[83]));
 sg13g2_buf_1 _1287_ (.A(net124),
    .X(results[84]));
 sg13g2_buf_1 _1288_ (.A(net125),
    .X(results[85]));
 sg13g2_buf_1 _1289_ (.A(net126),
    .X(results[86]));
 sg13g2_buf_1 _1290_ (.A(net127),
    .X(results[87]));
 sg13g2_buf_1 _1291_ (.A(net128),
    .X(results[88]));
 sg13g2_buf_1 _1292_ (.A(net129),
    .X(results[89]));
 sg13g2_buf_1 _1293_ (.A(net130),
    .X(results[90]));
 sg13g2_buf_1 _1294_ (.A(net131),
    .X(results[91]));
 sg13g2_buf_1 _1295_ (.A(net132),
    .X(results[92]));
 sg13g2_buf_1 _1296_ (.A(net133),
    .X(results[93]));
 sg13g2_buf_1 _1297_ (.A(net134),
    .X(results[94]));
 sg13g2_buf_1 _1298_ (.A(net135),
    .X(results[95]));
 sg13g2_buf_1 _1299_ (.A(net136),
    .X(results[96]));
 sg13g2_buf_1 _1300_ (.A(net137),
    .X(results[97]));
 sg13g2_buf_1 _1301_ (.A(net138),
    .X(results[98]));
 sg13g2_buf_1 _1302_ (.A(net139),
    .X(results[99]));
 sg13g2_buf_1 _1303_ (.A(net140),
    .X(results[100]));
 sg13g2_buf_1 _1304_ (.A(net141),
    .X(results[101]));
 sg13g2_buf_1 _1305_ (.A(net142),
    .X(results[102]));
 sg13g2_buf_1 _1306_ (.A(net143),
    .X(results[103]));
 sg13g2_buf_1 _1307_ (.A(net144),
    .X(results[104]));
 sg13g2_buf_1 _1308_ (.A(net145),
    .X(results[105]));
 sg13g2_buf_1 _1309_ (.A(net146),
    .X(results[106]));
 sg13g2_buf_1 _1310_ (.A(net147),
    .X(results[107]));
 sg13g2_buf_1 _1311_ (.A(net148),
    .X(results[112]));
 sg13g2_buf_1 _1312_ (.A(net149),
    .X(results[113]));
 sg13g2_buf_1 _1313_ (.A(net150),
    .X(results[114]));
 sg13g2_buf_1 _1314_ (.A(net151),
    .X(results[115]));
 sg13g2_buf_1 _1315_ (.A(net152),
    .X(results[116]));
 sg13g2_buf_1 _1316_ (.A(net153),
    .X(results[117]));
 sg13g2_buf_1 _1317_ (.A(net154),
    .X(results[118]));
 sg13g2_buf_1 _1318_ (.A(net155),
    .X(results[119]));
 sg13g2_buf_1 _1319_ (.A(net156),
    .X(results[120]));
 sg13g2_buf_1 _1320_ (.A(net157),
    .X(results[121]));
 sg13g2_buf_1 _1321_ (.A(net158),
    .X(results[122]));
 sg13g2_buf_1 _1322_ (.A(net159),
    .X(results[123]));
 sg13g2_buf_1 _1323_ (.A(net160),
    .X(results[124]));
 sg13g2_buf_1 _1324_ (.A(net161),
    .X(results[125]));
 sg13g2_buf_1 _1325_ (.A(net162),
    .X(results[126]));
 sg13g2_buf_1 _1326_ (.A(net163),
    .X(results[127]));
 sg13g2_dfrbp_1 \genblk1[0].pipe.counter[0]$_SDFFE_PP0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net164),
    .D(_0023_),
    .Q_N(_0636_),
    .Q(\genblk1[0].pipe.counter[0] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.counter[1]$_SDFFE_PP0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net165),
    .D(_0024_),
    .Q_N(_0635_),
    .Q(\genblk1[0].pipe.counter[1] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.counter[2]$_SDFFE_PP0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net166),
    .D(_0025_),
    .Q_N(_0634_),
    .Q(\genblk1[0].pipe.counter[2] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.counter[3]$_SDFFE_PP0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net167),
    .D(_0026_),
    .Q_N(_0633_),
    .Q(\genblk1[0].pipe.counter[3] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.counter[4]$_SDFFE_PP0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net168),
    .D(_0027_),
    .Q_N(_0632_),
    .Q(\genblk1[0].pipe.counter[4] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.result[12]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net169),
    .D(_0028_),
    .Q_N(_0631_),
    .Q(net39));
 sg13g2_dfrbp_1 \genblk1[0].pipe.result[13]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net170),
    .D(_0029_),
    .Q_N(_0630_),
    .Q(net40));
 sg13g2_dfrbp_1 \genblk1[0].pipe.result[14]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net171),
    .D(_0030_),
    .Q_N(_0629_),
    .Q(net41));
 sg13g2_dfrbp_1 \genblk1[0].pipe.result[15]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net172),
    .D(_0031_),
    .Q_N(_0637_),
    .Q(net42));
 sg13g2_dfrbp_1 \genblk1[0].pipe.state[0]$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net173),
    .D(_0000_),
    .Q_N(_0638_),
    .Q(\genblk1[0].pipe.state[0] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.state[1]$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net174),
    .D(_0001_),
    .Q_N(_0017_),
    .Q(\genblk1[0].pipe.state[1] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[24]$_SDFFE_PP0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net175),
    .D(_0032_),
    .Q_N(_0628_),
    .Q(\genblk1[0].pipe.eps[0][24] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[25]$_SDFFE_PP0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net176),
    .D(_0033_),
    .Q_N(_0627_),
    .Q(\genblk1[0].pipe.eps[0][25] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[26]$_SDFFE_PP0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net177),
    .D(_0034_),
    .Q_N(_0626_),
    .Q(\genblk1[0].pipe.eps[0][26] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[27]$_SDFFE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net178),
    .D(_0035_),
    .Q_N(_0008_),
    .Q(\genblk1[0].pipe.eps[0][27] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[28]$_SDFFE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net179),
    .D(_0036_),
    .Q_N(_0625_),
    .Q(\genblk1[0].pipe.eps[0][28] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[29]$_SDFFE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net180),
    .D(_0037_),
    .Q_N(_0013_),
    .Q(\genblk1[0].pipe.eps[0][29] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[30]$_SDFFE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net181),
    .D(_0038_),
    .Q_N(_0624_),
    .Q(\genblk1[0].pipe.eps[0][30] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.this_query[31]$_SDFFE_PP0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net182),
    .D(_0039_),
    .Q_N(_0011_),
    .Q(\genblk1[0].pipe.eps[0][31] ));
 sg13g2_dfrbp_1 \genblk1[0].pipe.valid$_SDFFE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net183),
    .D(_0040_),
    .Q_N(_0623_),
    .Q(\genblk1[0].pipe.valid ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.counter[0]$_SDFFE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net184),
    .D(_0041_),
    .Q_N(_0622_),
    .Q(\genblk1[1].pipe.counter[0] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.counter[1]$_SDFFE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net185),
    .D(_0042_),
    .Q_N(_0621_),
    .Q(\genblk1[1].pipe.counter[1] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.counter[2]$_SDFFE_PP0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net186),
    .D(_0043_),
    .Q_N(_0620_),
    .Q(\genblk1[1].pipe.counter[2] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.counter[3]$_SDFFE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net187),
    .D(_0044_),
    .Q_N(_0619_),
    .Q(\genblk1[1].pipe.counter[3] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.counter[4]$_SDFFE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net188),
    .D(_0045_),
    .Q_N(_0618_),
    .Q(\genblk1[1].pipe.counter[4] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.result[12]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net189),
    .D(_0046_),
    .Q_N(_0617_),
    .Q(net43));
 sg13g2_dfrbp_1 \genblk1[1].pipe.result[13]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net190),
    .D(_0047_),
    .Q_N(_0616_),
    .Q(net44));
 sg13g2_dfrbp_1 \genblk1[1].pipe.result[14]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net191),
    .D(_0048_),
    .Q_N(_0615_),
    .Q(net45));
 sg13g2_dfrbp_1 \genblk1[1].pipe.result[15]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net192),
    .D(_0049_),
    .Q_N(_0639_),
    .Q(net46));
 sg13g2_dfrbp_1 \genblk1[1].pipe.state[0]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net193),
    .D(_0002_),
    .Q_N(_0640_),
    .Q(\genblk1[1].pipe.state[0] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.state[1]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net194),
    .D(_0003_),
    .Q_N(_0019_),
    .Q(\genblk1[1].pipe.state[1] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[24]$_SDFFE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net195),
    .D(_0050_),
    .Q_N(_0614_),
    .Q(\genblk1[1].pipe.eps[0][24] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[25]$_SDFFE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net196),
    .D(_0051_),
    .Q_N(_0613_),
    .Q(\genblk1[1].pipe.eps[0][25] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[26]$_SDFFE_PP0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net197),
    .D(_0052_),
    .Q_N(_0612_),
    .Q(\genblk1[1].pipe.eps[0][26] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[27]$_SDFFE_PP0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net198),
    .D(_0053_),
    .Q_N(_0022_),
    .Q(\genblk1[1].pipe.eps[0][27] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[28]$_SDFFE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net199),
    .D(_0054_),
    .Q_N(_0611_),
    .Q(\genblk1[1].pipe.eps[0][28] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[29]$_SDFFE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net200),
    .D(_0055_),
    .Q_N(_0021_),
    .Q(\genblk1[1].pipe.eps[0][29] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[30]$_SDFFE_PP0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net201),
    .D(_0056_),
    .Q_N(_0610_),
    .Q(\genblk1[1].pipe.eps[0][30] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.this_query[31]$_SDFFE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net202),
    .D(_0057_),
    .Q_N(_0020_),
    .Q(\genblk1[1].pipe.eps[0][31] ));
 sg13g2_dfrbp_1 \genblk1[1].pipe.valid$_SDFFE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net203),
    .D(_0058_),
    .Q_N(_0609_),
    .Q(\genblk1[1].pipe.valid ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.counter[0]$_SDFFE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net204),
    .D(_0059_),
    .Q_N(_0608_),
    .Q(\genblk1[2].pipe.counter[0] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.counter[1]$_SDFFE_PP0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net205),
    .D(_0060_),
    .Q_N(_0607_),
    .Q(\genblk1[2].pipe.counter[1] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.counter[2]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net206),
    .D(_0061_),
    .Q_N(_0606_),
    .Q(\genblk1[2].pipe.counter[2] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.counter[3]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net207),
    .D(_0062_),
    .Q_N(_0605_),
    .Q(\genblk1[2].pipe.counter[3] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.counter[4]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net208),
    .D(_0063_),
    .Q_N(_0604_),
    .Q(\genblk1[2].pipe.counter[4] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.result[12]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net209),
    .D(_0064_),
    .Q_N(_0603_),
    .Q(net47));
 sg13g2_dfrbp_1 \genblk1[2].pipe.result[13]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net210),
    .D(_0065_),
    .Q_N(_0602_),
    .Q(net48));
 sg13g2_dfrbp_1 \genblk1[2].pipe.result[14]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net211),
    .D(_0066_),
    .Q_N(_0601_),
    .Q(net49));
 sg13g2_dfrbp_1 \genblk1[2].pipe.result[15]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net212),
    .D(_0067_),
    .Q_N(_0641_),
    .Q(net50));
 sg13g2_dfrbp_1 \genblk1[2].pipe.state[0]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net213),
    .D(_0004_),
    .Q_N(_0642_),
    .Q(\genblk1[2].pipe.state[0] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.state[1]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net214),
    .D(_0005_),
    .Q_N(_0009_),
    .Q(\genblk1[2].pipe.state[1] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[24]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net215),
    .D(_0068_),
    .Q_N(_0600_),
    .Q(\genblk1[2].pipe.eps[0][24] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[25]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net216),
    .D(_0069_),
    .Q_N(_0599_),
    .Q(\genblk1[2].pipe.eps[0][25] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[26]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net217),
    .D(_0070_),
    .Q_N(_0598_),
    .Q(\genblk1[2].pipe.eps[0][26] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[27]$_SDFFE_PP0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net218),
    .D(_0071_),
    .Q_N(_0018_),
    .Q(\genblk1[2].pipe.eps[0][27] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[28]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net219),
    .D(_0072_),
    .Q_N(_0597_),
    .Q(\genblk1[2].pipe.eps[0][28] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[29]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net220),
    .D(_0073_),
    .Q_N(_0016_),
    .Q(\genblk1[2].pipe.eps[0][29] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[30]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net221),
    .D(_0074_),
    .Q_N(_0596_),
    .Q(\genblk1[2].pipe.eps[0][30] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.this_query[31]$_SDFFE_PP0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net222),
    .D(_0075_),
    .Q_N(_0012_),
    .Q(\genblk1[2].pipe.eps[0][31] ));
 sg13g2_dfrbp_1 \genblk1[2].pipe.valid$_SDFFE_PP0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net223),
    .D(_0076_),
    .Q_N(_0595_),
    .Q(\genblk1[2].pipe.valid ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.counter[0]$_SDFFE_PP0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net224),
    .D(_0077_),
    .Q_N(_0594_),
    .Q(\genblk1[3].pipe.counter[0] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.counter[1]$_SDFFE_PP0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net225),
    .D(_0078_),
    .Q_N(_0593_),
    .Q(\genblk1[3].pipe.counter[1] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.counter[2]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net226),
    .D(_0079_),
    .Q_N(_0592_),
    .Q(\genblk1[3].pipe.counter[2] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.counter[3]$_SDFFE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net227),
    .D(_0080_),
    .Q_N(_0591_),
    .Q(\genblk1[3].pipe.counter[3] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.counter[4]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net228),
    .D(_0081_),
    .Q_N(_0590_),
    .Q(\genblk1[3].pipe.counter[4] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.result[12]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net229),
    .D(_0082_),
    .Q_N(_0589_),
    .Q(net35));
 sg13g2_dfrbp_1 \genblk1[3].pipe.result[13]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net230),
    .D(_0083_),
    .Q_N(_0588_),
    .Q(net36));
 sg13g2_dfrbp_1 \genblk1[3].pipe.result[14]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net231),
    .D(_0084_),
    .Q_N(_0587_),
    .Q(net37));
 sg13g2_dfrbp_1 \genblk1[3].pipe.result[15]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net232),
    .D(_0085_),
    .Q_N(_0643_),
    .Q(net38));
 sg13g2_dfrbp_1 \genblk1[3].pipe.state[0]$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net233),
    .D(_0006_),
    .Q_N(_0644_),
    .Q(\genblk1[3].pipe.state[0] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.state[1]$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net234),
    .D(_0007_),
    .Q_N(_0586_),
    .Q(\genblk1[3].pipe.state[1] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[24]$_SDFFE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net235),
    .D(_0086_),
    .Q_N(_0585_),
    .Q(\genblk1[3].pipe.eps[0][24] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[25]$_SDFFE_PP0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net236),
    .D(_0087_),
    .Q_N(_0584_),
    .Q(\genblk1[3].pipe.eps[0][25] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[26]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net237),
    .D(_0088_),
    .Q_N(_0583_),
    .Q(\genblk1[3].pipe.eps[0][26] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[27]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net238),
    .D(_0089_),
    .Q_N(_0010_),
    .Q(\genblk1[3].pipe.eps[0][27] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[28]$_SDFFE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net239),
    .D(_0090_),
    .Q_N(_0582_),
    .Q(\genblk1[3].pipe.eps[0][28] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[29]$_SDFFE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net240),
    .D(_0091_),
    .Q_N(_0014_),
    .Q(\genblk1[3].pipe.eps[0][29] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[30]$_SDFFE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net277),
    .D(_0092_),
    .Q_N(_0581_),
    .Q(\genblk1[3].pipe.eps[0][30] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.this_query[31]$_SDFFE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net278),
    .D(_0093_),
    .Q_N(_0015_),
    .Q(\genblk1[3].pipe.eps[0][31] ));
 sg13g2_dfrbp_1 \genblk1[3].pipe.valid$_SDFFE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net279),
    .D(_0094_),
    .Q_N(_0580_),
    .Q(\genblk1[3].pipe.valid ));
 sg13g2_tielo _1217__3 (.L_LO(net54));
 sg13g2_tielo _1223__9 (.L_LO(net60));
 sg13g2_buf_4 place241 (.X(net241),
    .A(_0167_));
 sg13g2_tielo _1219__5 (.L_LO(net56));
 sg13g2_tielo asqrt_top_1 (.L_LO(net52));
 sg13g2_tielo _1224__10 (.L_LO(net61));
 sg13g2_tielo _1227__13 (.L_LO(net64));
 sg13g2_buf_4 place244 (.X(net244),
    .A(_0538_));
 sg13g2_buf_4 place245 (.X(net245),
    .A(_0170_));
 sg13g2_buf_4 place270 (.X(net270),
    .A(net34));
 sg13g2_buf_4 place271 (.X(net271),
    .A(net270));
 sg13g2_tielo _1228__14 (.L_LO(net65));
 sg13g2_tielo _1229__15 (.L_LO(net66));
 sg13g2_tielo _1230__16 (.L_LO(net67));
 sg13g2_tielo _1231__17 (.L_LO(net68));
 sg13g2_tielo _1232__18 (.L_LO(net69));
 sg13g2_tielo _1233__19 (.L_LO(net70));
 sg13g2_tielo _1234__20 (.L_LO(net71));
 sg13g2_tielo _1235__21 (.L_LO(net72));
 sg13g2_tielo _1236__22 (.L_LO(net73));
 sg13g2_tielo _1237__23 (.L_LO(net74));
 sg13g2_tielo _1238__24 (.L_LO(net75));
 sg13g2_tielo _1239__25 (.L_LO(net76));
 sg13g2_tielo _1240__26 (.L_LO(net77));
 sg13g2_tielo _1241__27 (.L_LO(net78));
 sg13g2_tielo _1242__28 (.L_LO(net79));
 sg13g2_tielo _1243__29 (.L_LO(net80));
 sg13g2_tielo _1244__30 (.L_LO(net81));
 sg13g2_tielo _1245__31 (.L_LO(net82));
 sg13g2_tielo _1246__32 (.L_LO(net83));
 sg13g2_tielo _1247__33 (.L_LO(net84));
 sg13g2_tielo _1248__34 (.L_LO(net85));
 sg13g2_tielo _1249__35 (.L_LO(net86));
 sg13g2_tielo _1250__36 (.L_LO(net87));
 sg13g2_tielo _1251__37 (.L_LO(net88));
 sg13g2_tielo _1252__38 (.L_LO(net89));
 sg13g2_tielo _1253__39 (.L_LO(net90));
 sg13g2_tielo _1254__40 (.L_LO(net91));
 sg13g2_tielo _1255__41 (.L_LO(net92));
 sg13g2_tielo _1256__42 (.L_LO(net93));
 sg13g2_tielo _1257__43 (.L_LO(net94));
 sg13g2_tielo _1258__44 (.L_LO(net95));
 sg13g2_tielo _1259__45 (.L_LO(net96));
 sg13g2_tielo _1260__46 (.L_LO(net97));
 sg13g2_tielo _1261__47 (.L_LO(net98));
 sg13g2_tielo _1262__48 (.L_LO(net99));
 sg13g2_tielo _1263__49 (.L_LO(net100));
 sg13g2_tielo _1264__50 (.L_LO(net101));
 sg13g2_tielo _1265__51 (.L_LO(net102));
 sg13g2_tielo _1266__52 (.L_LO(net103));
 sg13g2_tielo _1267__53 (.L_LO(net104));
 sg13g2_tielo _1268__54 (.L_LO(net105));
 sg13g2_tielo _1269__55 (.L_LO(net106));
 sg13g2_tielo _1270__56 (.L_LO(net107));
 sg13g2_tielo _1271__57 (.L_LO(net108));
 sg13g2_tielo _1272__58 (.L_LO(net109));
 sg13g2_tielo _1273__59 (.L_LO(net110));
 sg13g2_tielo _1274__60 (.L_LO(net111));
 sg13g2_tielo _1275__61 (.L_LO(net112));
 sg13g2_tielo _1276__62 (.L_LO(net113));
 sg13g2_tielo _1277__63 (.L_LO(net114));
 sg13g2_tielo _1278__64 (.L_LO(net115));
 sg13g2_tielo _1279__65 (.L_LO(net116));
 sg13g2_tielo _1280__66 (.L_LO(net117));
 sg13g2_tielo _1281__67 (.L_LO(net118));
 sg13g2_tielo _1282__68 (.L_LO(net119));
 sg13g2_tielo _1283__69 (.L_LO(net120));
 sg13g2_tielo _1284__70 (.L_LO(net121));
 sg13g2_tielo _1285__71 (.L_LO(net122));
 sg13g2_tielo _1286__72 (.L_LO(net123));
 sg13g2_tielo _1287__73 (.L_LO(net124));
 sg13g2_tielo _1288__74 (.L_LO(net125));
 sg13g2_tielo _1289__75 (.L_LO(net126));
 sg13g2_tielo _1290__76 (.L_LO(net127));
 sg13g2_tielo _1291__77 (.L_LO(net128));
 sg13g2_tielo _1292__78 (.L_LO(net129));
 sg13g2_tielo _1293__79 (.L_LO(net130));
 sg13g2_tielo _1294__80 (.L_LO(net131));
 sg13g2_tielo _1295__81 (.L_LO(net132));
 sg13g2_tielo _1296__82 (.L_LO(net133));
 sg13g2_tielo _1297__83 (.L_LO(net134));
 sg13g2_tielo _1298__84 (.L_LO(net135));
 sg13g2_tielo _1299__85 (.L_LO(net136));
 sg13g2_tielo _1300__86 (.L_LO(net137));
 sg13g2_tielo _1301__87 (.L_LO(net138));
 sg13g2_tielo _1302__88 (.L_LO(net139));
 sg13g2_tielo _1303__89 (.L_LO(net140));
 sg13g2_tielo _1304__90 (.L_LO(net141));
 sg13g2_tielo _1305__91 (.L_LO(net142));
 sg13g2_tielo _1306__92 (.L_LO(net143));
 sg13g2_tielo _1307__93 (.L_LO(net144));
 sg13g2_tielo _1308__94 (.L_LO(net145));
 sg13g2_tielo _1309__95 (.L_LO(net146));
 sg13g2_tielo _1310__96 (.L_LO(net147));
 sg13g2_tielo _1311__97 (.L_LO(net148));
 sg13g2_tielo _1312__98 (.L_LO(net149));
 sg13g2_tielo _1313__99 (.L_LO(net150));
 sg13g2_tielo _1314__100 (.L_LO(net151));
 sg13g2_tielo _1315__101 (.L_LO(net152));
 sg13g2_tielo _1316__102 (.L_LO(net153));
 sg13g2_tielo _1317__103 (.L_LO(net154));
 sg13g2_tielo _1318__104 (.L_LO(net155));
 sg13g2_tielo _1319__105 (.L_LO(net156));
 sg13g2_tielo _1320__106 (.L_LO(net157));
 sg13g2_tielo _1321__107 (.L_LO(net158));
 sg13g2_tielo _1322__108 (.L_LO(net159));
 sg13g2_tielo _1323__109 (.L_LO(net160));
 sg13g2_tielo _1324__110 (.L_LO(net161));
 sg13g2_tielo _1325__111 (.L_LO(net162));
 sg13g2_tielo _1326__112 (.L_LO(net163));
 sg13g2_tiehi \genblk1[0].pipe.counter[1]$_SDFFE_PP0P__114  (.L_HI(net165));
 sg13g2_tiehi \genblk1[0].pipe.counter[2]$_SDFFE_PP0P__115  (.L_HI(net166));
 sg13g2_tiehi \genblk1[0].pipe.counter[3]$_SDFFE_PP0P__116  (.L_HI(net167));
 sg13g2_tiehi \genblk1[0].pipe.counter[4]$_SDFFE_PP0P__117  (.L_HI(net168));
 sg13g2_tiehi \genblk1[0].pipe.result[12]$_DFFE_PP__118  (.L_HI(net169));
 sg13g2_tiehi \genblk1[0].pipe.result[13]$_DFFE_PP__119  (.L_HI(net170));
 sg13g2_tiehi \genblk1[0].pipe.result[14]$_DFFE_PP__120  (.L_HI(net171));
 sg13g2_tiehi \genblk1[0].pipe.result[15]$_DFFE_PP__121  (.L_HI(net172));
 sg13g2_tiehi \genblk1[0].pipe.state[0]$_DFF_P__122  (.L_HI(net173));
 sg13g2_tiehi \genblk1[0].pipe.state[1]$_DFF_P__123  (.L_HI(net174));
 sg13g2_tiehi \genblk1[0].pipe.this_query[24]$_SDFFE_PP0P__124  (.L_HI(net175));
 sg13g2_tiehi \genblk1[0].pipe.this_query[25]$_SDFFE_PP0P__125  (.L_HI(net176));
 sg13g2_tiehi \genblk1[0].pipe.this_query[26]$_SDFFE_PP0P__126  (.L_HI(net177));
 sg13g2_tiehi \genblk1[0].pipe.this_query[27]$_SDFFE_PP0P__127  (.L_HI(net178));
 sg13g2_tiehi \genblk1[0].pipe.this_query[28]$_SDFFE_PP0P__128  (.L_HI(net179));
 sg13g2_tiehi \genblk1[0].pipe.this_query[29]$_SDFFE_PP0P__129  (.L_HI(net180));
 sg13g2_tiehi \genblk1[0].pipe.this_query[30]$_SDFFE_PP0P__130  (.L_HI(net181));
 sg13g2_tiehi \genblk1[0].pipe.this_query[31]$_SDFFE_PP0P__131  (.L_HI(net182));
 sg13g2_tiehi \genblk1[0].pipe.valid$_SDFFE_PP0P__132  (.L_HI(net183));
 sg13g2_tiehi \genblk1[1].pipe.counter[0]$_SDFFE_PP0P__133  (.L_HI(net184));
 sg13g2_tiehi \genblk1[1].pipe.counter[1]$_SDFFE_PP0P__134  (.L_HI(net185));
 sg13g2_tiehi \genblk1[1].pipe.counter[2]$_SDFFE_PP0P__135  (.L_HI(net186));
 sg13g2_tiehi \genblk1[1].pipe.counter[3]$_SDFFE_PP0P__136  (.L_HI(net187));
 sg13g2_tiehi \genblk1[1].pipe.counter[4]$_SDFFE_PP0P__137  (.L_HI(net188));
 sg13g2_tiehi \genblk1[1].pipe.result[12]$_DFFE_PP__138  (.L_HI(net189));
 sg13g2_tiehi \genblk1[1].pipe.result[13]$_DFFE_PP__139  (.L_HI(net190));
 sg13g2_tiehi \genblk1[1].pipe.result[14]$_DFFE_PP__140  (.L_HI(net191));
 sg13g2_tiehi \genblk1[1].pipe.result[15]$_DFFE_PP__141  (.L_HI(net192));
 sg13g2_tiehi \genblk1[1].pipe.state[0]$_DFF_P__142  (.L_HI(net193));
 sg13g2_tiehi \genblk1[1].pipe.state[1]$_DFF_P__143  (.L_HI(net194));
 sg13g2_tiehi \genblk1[1].pipe.this_query[24]$_SDFFE_PP0P__144  (.L_HI(net195));
 sg13g2_tiehi \genblk1[1].pipe.this_query[25]$_SDFFE_PP0P__145  (.L_HI(net196));
 sg13g2_tiehi \genblk1[1].pipe.this_query[26]$_SDFFE_PP0P__146  (.L_HI(net197));
 sg13g2_tiehi \genblk1[1].pipe.this_query[27]$_SDFFE_PP0P__147  (.L_HI(net198));
 sg13g2_tiehi \genblk1[1].pipe.this_query[28]$_SDFFE_PP0P__148  (.L_HI(net199));
 sg13g2_tiehi \genblk1[1].pipe.this_query[29]$_SDFFE_PP0P__149  (.L_HI(net200));
 sg13g2_tiehi \genblk1[1].pipe.this_query[30]$_SDFFE_PP0P__150  (.L_HI(net201));
 sg13g2_tiehi \genblk1[1].pipe.this_query[31]$_SDFFE_PP0P__151  (.L_HI(net202));
 sg13g2_tiehi \genblk1[1].pipe.valid$_SDFFE_PP0P__152  (.L_HI(net203));
 sg13g2_tiehi \genblk1[2].pipe.counter[0]$_SDFFE_PP0P__153  (.L_HI(net204));
 sg13g2_tiehi \genblk1[2].pipe.counter[1]$_SDFFE_PP0P__154  (.L_HI(net205));
 sg13g2_tiehi \genblk1[2].pipe.counter[2]$_SDFFE_PP0P__155  (.L_HI(net206));
 sg13g2_tiehi \genblk1[2].pipe.counter[3]$_SDFFE_PP0P__156  (.L_HI(net207));
 sg13g2_tiehi \genblk1[2].pipe.counter[4]$_SDFFE_PP0P__157  (.L_HI(net208));
 sg13g2_tiehi \genblk1[2].pipe.result[12]$_DFFE_PP__158  (.L_HI(net209));
 sg13g2_tiehi \genblk1[2].pipe.result[13]$_DFFE_PP__159  (.L_HI(net210));
 sg13g2_tiehi \genblk1[2].pipe.result[14]$_DFFE_PP__160  (.L_HI(net211));
 sg13g2_tiehi \genblk1[2].pipe.result[15]$_DFFE_PP__161  (.L_HI(net212));
 sg13g2_tiehi \genblk1[2].pipe.state[0]$_DFF_P__162  (.L_HI(net213));
 sg13g2_tiehi \genblk1[2].pipe.state[1]$_DFF_P__163  (.L_HI(net214));
 sg13g2_tiehi \genblk1[2].pipe.this_query[24]$_SDFFE_PP0P__164  (.L_HI(net215));
 sg13g2_tiehi \genblk1[2].pipe.this_query[25]$_SDFFE_PP0P__165  (.L_HI(net216));
 sg13g2_tiehi \genblk1[2].pipe.this_query[26]$_SDFFE_PP0P__166  (.L_HI(net217));
 sg13g2_tiehi \genblk1[2].pipe.this_query[27]$_SDFFE_PP0P__167  (.L_HI(net218));
 sg13g2_tiehi \genblk1[2].pipe.this_query[28]$_SDFFE_PP0P__168  (.L_HI(net219));
 sg13g2_tiehi \genblk1[2].pipe.this_query[29]$_SDFFE_PP0P__169  (.L_HI(net220));
 sg13g2_tiehi \genblk1[2].pipe.this_query[30]$_SDFFE_PP0P__170  (.L_HI(net221));
 sg13g2_tiehi \genblk1[2].pipe.this_query[31]$_SDFFE_PP0P__171  (.L_HI(net222));
 sg13g2_tiehi \genblk1[2].pipe.valid$_SDFFE_PP0P__172  (.L_HI(net223));
 sg13g2_tiehi \genblk1[3].pipe.counter[0]$_SDFFE_PP0P__173  (.L_HI(net224));
 sg13g2_tiehi \genblk1[3].pipe.counter[1]$_SDFFE_PP0P__174  (.L_HI(net225));
 sg13g2_tiehi \genblk1[3].pipe.counter[2]$_SDFFE_PP0P__175  (.L_HI(net226));
 sg13g2_tiehi \genblk1[3].pipe.counter[3]$_SDFFE_PP0P__176  (.L_HI(net227));
 sg13g2_tiehi \genblk1[3].pipe.counter[4]$_SDFFE_PP0P__177  (.L_HI(net228));
 sg13g2_tiehi \genblk1[3].pipe.result[12]$_DFFE_PP__178  (.L_HI(net229));
 sg13g2_tiehi \genblk1[3].pipe.result[13]$_DFFE_PP__179  (.L_HI(net230));
 sg13g2_tiehi \genblk1[3].pipe.result[14]$_DFFE_PP__180  (.L_HI(net231));
 sg13g2_tiehi \genblk1[3].pipe.result[15]$_DFFE_PP__181  (.L_HI(net232));
 sg13g2_tiehi \genblk1[3].pipe.state[0]$_DFF_P__182  (.L_HI(net233));
 sg13g2_tiehi \genblk1[3].pipe.state[1]$_DFF_P__183  (.L_HI(net234));
 sg13g2_tiehi \genblk1[3].pipe.this_query[24]$_SDFFE_PP0P__184  (.L_HI(net235));
 sg13g2_tiehi \genblk1[3].pipe.this_query[25]$_SDFFE_PP0P__185  (.L_HI(net236));
 sg13g2_tiehi \genblk1[3].pipe.this_query[26]$_SDFFE_PP0P__186  (.L_HI(net237));
 sg13g2_tiehi \genblk1[3].pipe.this_query[27]$_SDFFE_PP0P__187  (.L_HI(net238));
 sg13g2_tiehi \genblk1[3].pipe.this_query[28]$_SDFFE_PP0P__188  (.L_HI(net239));
 sg13g2_tiehi \genblk1[3].pipe.this_query[29]$_SDFFE_PP0P__189  (.L_HI(net240));
 sg13g2_tiehi \genblk1[3].pipe.this_query[30]$_SDFFE_PP0P__190  (.L_HI(net277));
 sg13g2_tiehi \genblk1[3].pipe.this_query[31]$_SDFFE_PP0P__191  (.L_HI(net278));
 sg13g2_tiehi \genblk1[3].pipe.valid$_SDFFE_PP0P__192  (.L_HI(net279));
 sg13g2_buf_16 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1 (.A(queries[124]));
 sg13g2_antennanp ANTENNA_2 (.A(queries[125]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_fill_2 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_4 FILLER_0_326 ();
 sg13g2_fill_1 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_fill_2 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_166 ();
 sg13g2_fill_1 FILLER_1_196 ();
 sg13g2_decap_4 FILLER_1_202 ();
 sg13g2_decap_8 FILLER_1_247 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_decap_8 FILLER_1_261 ();
 sg13g2_decap_8 FILLER_1_268 ();
 sg13g2_decap_8 FILLER_1_275 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_fill_2 FILLER_2_123 ();
 sg13g2_fill_1 FILLER_2_125 ();
 sg13g2_decap_4 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_165 ();
 sg13g2_decap_4 FILLER_2_222 ();
 sg13g2_fill_1 FILLER_2_229 ();
 sg13g2_fill_2 FILLER_2_235 ();
 sg13g2_fill_1 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_248 ();
 sg13g2_decap_8 FILLER_2_255 ();
 sg13g2_decap_8 FILLER_2_262 ();
 sg13g2_decap_8 FILLER_2_269 ();
 sg13g2_decap_8 FILLER_2_276 ();
 sg13g2_decap_8 FILLER_2_283 ();
 sg13g2_decap_8 FILLER_2_290 ();
 sg13g2_decap_8 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_4 FILLER_2_325 ();
 sg13g2_fill_2 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_4 FILLER_3_84 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_115 ();
 sg13g2_decap_4 FILLER_3_122 ();
 sg13g2_fill_1 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_fill_2 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_152 ();
 sg13g2_decap_4 FILLER_3_167 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_1 FILLER_3_191 ();
 sg13g2_fill_2 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_251 ();
 sg13g2_decap_8 FILLER_3_258 ();
 sg13g2_decap_8 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_279 ();
 sg13g2_decap_8 FILLER_3_286 ();
 sg13g2_decap_8 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_300 ();
 sg13g2_decap_8 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_321 ();
 sg13g2_fill_2 FILLER_3_328 ();
 sg13g2_fill_1 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_4 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_fill_2 FILLER_4_84 ();
 sg13g2_fill_1 FILLER_4_86 ();
 sg13g2_decap_4 FILLER_4_92 ();
 sg13g2_fill_2 FILLER_4_96 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_4 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_131 ();
 sg13g2_fill_2 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_145 ();
 sg13g2_decap_8 FILLER_4_152 ();
 sg13g2_decap_8 FILLER_4_159 ();
 sg13g2_decap_8 FILLER_4_166 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_fill_2 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_232 ();
 sg13g2_fill_1 FILLER_4_234 ();
 sg13g2_decap_8 FILLER_4_244 ();
 sg13g2_decap_8 FILLER_4_251 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_decap_8 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_272 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_decap_8 FILLER_4_314 ();
 sg13g2_decap_8 FILLER_4_321 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_fill_2 FILLER_5_42 ();
 sg13g2_fill_1 FILLER_5_83 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_4 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_180 ();
 sg13g2_decap_8 FILLER_5_187 ();
 sg13g2_decap_8 FILLER_5_194 ();
 sg13g2_decap_8 FILLER_5_201 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_4 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_decap_8 FILLER_5_269 ();
 sg13g2_decap_8 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_4 FILLER_5_325 ();
 sg13g2_fill_2 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_115 ();
 sg13g2_fill_1 FILLER_6_122 ();
 sg13g2_fill_2 FILLER_6_127 ();
 sg13g2_fill_1 FILLER_6_129 ();
 sg13g2_decap_4 FILLER_6_160 ();
 sg13g2_fill_1 FILLER_6_169 ();
 sg13g2_decap_8 FILLER_6_209 ();
 sg13g2_decap_8 FILLER_6_216 ();
 sg13g2_decap_8 FILLER_6_223 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_4 FILLER_6_325 ();
 sg13g2_fill_2 FILLER_6_329 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_4 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_47 ();
 sg13g2_decap_8 FILLER_7_54 ();
 sg13g2_decap_8 FILLER_7_61 ();
 sg13g2_decap_4 FILLER_7_82 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_fill_2 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_4 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_9 ();
 sg13g2_decap_4 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_fill_1 FILLER_8_59 ();
 sg13g2_decap_4 FILLER_8_85 ();
 sg13g2_decap_4 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_150 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_219 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_fill_1 FILLER_8_237 ();
 sg13g2_fill_1 FILLER_8_248 ();
 sg13g2_fill_1 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_fill_1 FILLER_8_330 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_decap_4 FILLER_9_16 ();
 sg13g2_fill_2 FILLER_9_20 ();
 sg13g2_fill_1 FILLER_9_27 ();
 sg13g2_fill_1 FILLER_9_33 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_fill_2 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_89 ();
 sg13g2_fill_1 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_4 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_240 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_13 ();
 sg13g2_decap_4 FILLER_10_23 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_4 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_43 ();
 sg13g2_fill_2 FILLER_10_48 ();
 sg13g2_fill_2 FILLER_10_64 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_4 FILLER_10_81 ();
 sg13g2_fill_2 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_92 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_4 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_fill_1 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_4 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_4 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_45 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_71 ();
 sg13g2_decap_8 FILLER_11_86 ();
 sg13g2_decap_8 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_104 ();
 sg13g2_decap_8 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_125 ();
 sg13g2_decap_4 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_decap_4 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_151 ();
 sg13g2_fill_2 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_171 ();
 sg13g2_decap_8 FILLER_11_178 ();
 sg13g2_decap_8 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_decap_4 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_4 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_329 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_decap_4 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_26 ();
 sg13g2_decap_8 FILLER_12_33 ();
 sg13g2_decap_8 FILLER_12_40 ();
 sg13g2_fill_1 FILLER_12_47 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_54 ();
 sg13g2_decap_4 FILLER_12_89 ();
 sg13g2_decap_8 FILLER_12_104 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_fill_2 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_211 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_4 FILLER_12_326 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_33 ();
 sg13g2_decap_8 FILLER_13_40 ();
 sg13g2_fill_1 FILLER_13_47 ();
 sg13g2_decap_8 FILLER_13_89 ();
 sg13g2_decap_8 FILLER_13_96 ();
 sg13g2_decap_8 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_4 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_264 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_4 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_37 ();
 sg13g2_decap_8 FILLER_14_44 ();
 sg13g2_fill_1 FILLER_14_51 ();
 sg13g2_decap_8 FILLER_14_78 ();
 sg13g2_decap_4 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_89 ();
 sg13g2_decap_4 FILLER_14_94 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_fill_2 FILLER_14_132 ();
 sg13g2_decap_4 FILLER_14_139 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_decap_4 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_fill_2 FILLER_14_169 ();
 sg13g2_fill_1 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_31 ();
 sg13g2_decap_8 FILLER_15_38 ();
 sg13g2_decap_8 FILLER_15_45 ();
 sg13g2_decap_8 FILLER_15_52 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_75 ();
 sg13g2_fill_2 FILLER_15_82 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_4 FILLER_15_130 ();
 sg13g2_fill_2 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_4 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_181 ();
 sg13g2_decap_4 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_decap_4 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_decap_4 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_15 ();
 sg13g2_fill_2 FILLER_16_22 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_decap_8 FILLER_16_73 ();
 sg13g2_decap_8 FILLER_16_80 ();
 sg13g2_fill_1 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_4 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_4 FILLER_16_240 ();
 sg13g2_decap_4 FILLER_16_267 ();
 sg13g2_decap_4 FILLER_16_275 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_11 ();
 sg13g2_decap_4 FILLER_17_15 ();
 sg13g2_fill_1 FILLER_17_19 ();
 sg13g2_fill_1 FILLER_17_37 ();
 sg13g2_fill_1 FILLER_17_43 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_1 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_79 ();
 sg13g2_decap_4 FILLER_17_86 ();
 sg13g2_fill_1 FILLER_17_95 ();
 sg13g2_decap_4 FILLER_17_152 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_decap_4 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_4 FILLER_17_233 ();
 sg13g2_decap_4 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_249 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_decap_4 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_9 ();
 sg13g2_decap_8 FILLER_18_45 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_69 ();
 sg13g2_decap_8 FILLER_18_85 ();
 sg13g2_decap_8 FILLER_18_92 ();
 sg13g2_fill_2 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_decap_4 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_decap_4 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_32 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_fill_2 FILLER_19_50 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_4 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_4 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_4 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_40 ();
 sg13g2_fill_2 FILLER_20_47 ();
 sg13g2_fill_1 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_4 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_decap_4 FILLER_20_122 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_188 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_decap_4 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_23 ();
 sg13g2_decap_8 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_295 ();
 sg13g2_fill_1 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_decap_8 FILLER_22_61 ();
 sg13g2_decap_8 FILLER_22_68 ();
 sg13g2_fill_2 FILLER_22_101 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_4 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_56 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_decap_4 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_4 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_102 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_62 ();
 sg13g2_decap_8 FILLER_25_69 ();
 sg13g2_decap_4 FILLER_25_76 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_257 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_299 ();
 sg13g2_fill_2 FILLER_25_314 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_90 ();
 sg13g2_decap_4 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_109 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_4 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_8 FILLER_26_163 ();
 sg13g2_decap_8 FILLER_26_170 ();
 sg13g2_decap_8 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_decap_4 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_4 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_decap_4 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_4 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_decap_4 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_fill_2 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_decap_4 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_decap_4 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_4 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_4 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_decap_8 FILLER_29_117 ();
 sg13g2_decap_8 FILLER_29_124 ();
 sg13g2_decap_4 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_155 ();
 sg13g2_decap_4 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_166 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_194 ();
 sg13g2_decap_4 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_211 ();
 sg13g2_decap_4 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_4 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_157 ();
 sg13g2_decap_8 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_decap_4 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_8 FILLER_31_310 ();
 sg13g2_decap_4 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_decap_4 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_160 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_decap_4 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_230 ();
 sg13g2_decap_4 FILLER_32_236 ();
 sg13g2_decap_4 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_fill_1 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_64 ();
 sg13g2_decap_8 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_decap_8 FILLER_33_85 ();
 sg13g2_decap_8 FILLER_33_92 ();
 sg13g2_decap_8 FILLER_33_99 ();
 sg13g2_decap_4 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_4 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_decap_4 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_53 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_fill_2 FILLER_34_76 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_decap_4 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_150 ();
 sg13g2_decap_8 FILLER_35_157 ();
 sg13g2_decap_8 FILLER_35_164 ();
 sg13g2_decap_8 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_178 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_decap_8 FILLER_35_220 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_60 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_2 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_decap_4 FILLER_36_128 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_decap_4 FILLER_36_240 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_88 ();
 sg13g2_fill_2 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_decap_4 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_4 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_fill_1 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_decap_4 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_234 ();
 sg13g2_decap_4 FILLER_38_246 ();
 sg13g2_decap_4 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_decap_4 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_88 ();
 sg13g2_decap_4 FILLER_39_95 ();
 sg13g2_fill_2 FILLER_39_116 ();
 sg13g2_fill_1 FILLER_39_118 ();
 sg13g2_decap_4 FILLER_39_127 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_210 ();
 sg13g2_fill_1 FILLER_39_212 ();
 sg13g2_fill_1 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_238 ();
 sg13g2_fill_1 FILLER_39_247 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_fill_1 FILLER_39_287 ();
 sg13g2_fill_1 FILLER_39_292 ();
 sg13g2_fill_1 FILLER_39_305 ();
 sg13g2_fill_1 FILLER_39_330 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_236 ();
 sg13g2_fill_1 FILLER_40_241 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_282 ();
 sg13g2_fill_2 FILLER_40_291 ();
 sg13g2_fill_1 FILLER_40_293 ();
 sg13g2_fill_1 FILLER_40_326 ();
 assign results[0] = net52;
endmodule
